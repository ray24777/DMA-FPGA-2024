module axi_ahblite_top_45df1ab5d994#(
   parameter                    AL_US_AXI_ADDR_WIDTH = 32,      //Range: 32-64.
   parameter                    AL_US_AXI_DATA_WIDTH = 32,      //Range: 32,64.
   parameter                    AL_US_AXI_ID_WIDTH = 4,         //Range: 1-16.
   parameter                    AL_DS_AHB_ADDR_WIDTH = 32,      //Range: 32-64. !!AXI_ADDR_WIDTH = AHB_ADDR_WIDTH!!.
   parameter                    AL_DS_AHB_DATA_WIDTH = 32,      //Range: 32,64  !!AXI_DATA_WIDTH = AHB_DATA_WIDTH!!.
   parameter                    AL_SUPPORTS_NARROW_BURST = 1,   //Range: 0,1.   0:OFF  1:ON
   parameter                    AL_TIMEOUT_CYCLE = 16            //Range: 0,16,32,64,128,256.
)(
//Global signal
   input                              aclk,
   input                              aresetn,
//----------------AXI_Slave-------------------------
//AXI WADDR   
   input [AL_US_AXI_ID_WIDTH-1:0]     us_axi_awid,
   input [7:0]                        us_axi_awlen,
   input [2:0]                        us_axi_awsize,
   input [1:0]                        us_axi_awburst,
   input [3:0]                        us_axi_awcache,
   input [AL_US_AXI_ADDR_WIDTH-1:0]   us_axi_awaddr,
   input [2:0]                        us_axi_awprot,
   input                              us_axi_awvalid,
   output                             us_axi_awready,
   input                              us_axi_awlock,
//AXI WDATA
   input [AL_US_AXI_DATA_WIDTH-1:0]   us_axi_wdata,
   input [(AL_US_AXI_DATA_WIDTH/8)-1:0] us_axi_wstrb,
   input                              us_axi_wlast,
   input                              us_axi_wvalid,
   output                             us_axi_wready,
//AXI WRESP   
   output [AL_US_AXI_ID_WIDTH-1:0]    us_axi_bid,
   output [1:0]                       us_axi_bresp,
   output                             us_axi_bvalid,
   input                              us_axi_bready,
//AXI RADDR   
   input [AL_US_AXI_ID_WIDTH-1:0]     us_axi_arid,
   input [AL_US_AXI_ADDR_WIDTH-1:0]   us_axi_araddr,
   input [2:0]                        us_axi_arprot,
   input [3:0]                        us_axi_arcache,
   input                              us_axi_arvalid,
   input [7:0]                        us_axi_arlen,
   input [2:0]                        us_axi_arsize,
   input [1:0]                        us_axi_arburst,
   input                              us_axi_arlock,
   output                             us_axi_arready,
//AXI RDATA
   output [AL_US_AXI_ID_WIDTH-1:0]    us_axi_rid,
   output [AL_US_AXI_DATA_WIDTH-1:0]  us_axi_rdata,
   output [1:0]                       us_axi_rresp,
   output                             us_axi_rvalid,
   output                             us_axi_rlast,
   input                              us_axi_rready,
//-------------------AHB_Lite_Master----------------------  
   output [AL_DS_AHB_ADDR_WIDTH-1:0]  ds_ahb_haddr,
   output                             ds_ahb_hwrite,
   output [2:0]                       ds_ahb_hsize,
   output [2:0]                       ds_ahb_hburst,
   output [3:0]                       ds_ahb_hprot,
   output [1:0]                       ds_ahb_htrans,
   output                             ds_ahb_hmastlock,
   output [AL_DS_AHB_DATA_WIDTH-1:0]  ds_ahb_hwdata,
   
   input                              ds_ahb_hready,
   input [AL_DS_AHB_DATA_WIDTH-1:0]   ds_ahb_hrdata,
   input                              ds_ahb_hresp
    );
   `pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-009"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
m9qcOt5lHUz/F+lrpf6AiPTCWKXE3qqNfJG/HFNRiZ0nckVPx97nc4RMEMTbPAlf
9JGllIgoMFJ7ZH7Ezb7aOPNJkSQm4Bk5XljwMlN4C3xCMI0ALM9VstD55LiHiPF+
RlscFeoorMmSjhfzHHXPzK4LuaUOKjgOInTrRS6PuTI=
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
iGDe174QOvlGg6aywFQXo7uWAhN4/9k0obvYWOWGusqCpX9dMpkOLvV7wn9pURJJ
SVc/k6ZrdDNN54sV3nhuoebBnew1pJT7xrjeSzcFzxk5klM/XPFpyB0LuSobaLEt
AH29AJGazQi9huI94TG7Uid9Arrcpb8c8zYWSAU51rNwORcwx6yzeWBNnYzBaEIW
3Pdv72fMiZwPyCaHLc6l4VLbXh7eqhvCUUDZ6vVDVPZdRmqR04y3M3R8e1LIzaqU
WT1w8/ICWtGI1T1T5KAUprM9gvKBqTlxa/shvKs5Iou0UTuWvWaWHONuz5HY/E/i
WjSC4J10hdZZX/ROXMGQ9g==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
l0h7NRg/On5Dx1GbkkoiNzM4bC+6eT9ViAio4lpYNxma0uN6wih4hhZ6FxApwRvD
/2z+8eIPycdOWy0UQi8jO7G1vIsxHrh/drjoKGuNW/afFzmuH6+W8erpvHj6o1vc
P6gVW6u0emiyfnga4TCrq4yZyriMaa8UdwM5pNVqnog=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 89664)
`pragma protect data_block
cUizKmd7oPh2xiQZDVcoDVqsanb5dDH9RvYs+/vJOhm5Ztmkqx9+tZ1fJ2jNXBHK
7k7jyygaqObVD9ZZsR2+sXE8ZE6wzkKBW+4RSinmxj1yItqo6IZRPYx83tVpddY8
YjXbmb7kuC42N63P2e+hxgyHmjBg6U8EqJ0GslT6dsyx2fvt8qSJ8Ig4/vO6V9SA
tUvYuDnRrdDKkb4Sxaw9NsyPrre3NE74GnUzVXKcDnnwYBX3CwaYnaG08S1gknZj
Q9qJtK0G8tvF7c/b13T3T0A7Fz7yu9g5WFXF2KWBoNH8Lrcsr29WgfzBbOCs218e
oI95aWbfdCwO4G47rEG3LzJt+DNNFHxuJ1L7WuPSNopOcTjdtBlbxdyg39H9SdMQ
I2zBjedwA2h0HMgDZ/Y54jn6Cvi854vvQDbKNhdnvgQOCGnDc/NOTqyluwXuJV2n
yGJ3ymHvDHBTt11E/vITFxA444ykx/krHq9IERwJwOj5tzdbzAimg1p1LD0sFm4H
1u/Y3G9sKQiKwpZNaoDkBIrIGNfNUqRwMFfmnGWp/vJh4ggWuE8NnhiRWfv0jMhU
/KrGdA2cYpT4St5nkyY/ZXGFkoAZdZUEuvqbwKptL3V+7XqdQwyZdxVLUx9nv5Bi
pykQM59Mb4SWbs4AzeGvOvS/fi/YKkHcKwcp10VIfWNSIbxh6qALOF0I06gCOk68
ykm1NpMMTDjVysBI56x7IS64w/GPtwOpxJPNvfJGP3IlJNNG1y5ypNDOaWsYnnHi
/WHoXXB+7sKDzD7Gi0uYly+Cr99FZWB7ZTX+u1Uh0RE0tefM5YNWMWk5F5CHtKnb
e3VWbevAOhlfjM8zXITDde6R69+sl90Oct37vYHhWkX4/BR4iBgvhgmTnU6A8pRH
XgvzFufw99J0rnYvPqX+OycaKUTYX5dO7rc/BSNSH08RmmWWNh50Re12dkR6GVZV
H1YrtvVDWbCGBO+nTRQ9xU8OzW37W/qK2dxJxBpzXxHm/QrqOlxJXgzFx1eBn0aC
pjzb3BlXn/aBsmqwzOmOq8nJ//8M4iyZ7+4AN31MAA8lliZQebX3OGxM8CrQBEmY
U0FdOuxmBWI7FuFj385+iLdnlP6TruxxXQ6mfMPhF2pFUIt/yxcyYjFB1PXgtFpL
INy0rPqeM5kZjDgG+Gdlst87nz0jUjanYmiW5zo1r4jtkR86GcPBOtaRVjAuytC8
6sRw0T3l/jYhGZvnR3AxHPkWBKVdC1NsuKzmw8bKugCwgTXvR4fvnwXAY+XHiDt6
1PuBvl6O8rbBKYTnSHIZljtIIwDzUT59B9A5YlPzGW9TfsWUsT8UHddYbNAoikyn
Nn8j0JkqqyRaHTMIKdZSNq0N/bchEgfgeSosiq5OKkezZ5l9pkKCD7KctOFNk6kf
7HqAdwQS3EMY8r0KDhMUKf8sx6tFf460dshAinpSwugwWVuA1NMW2JYA3ej8p5jZ
PU0lhMkbNhCtldqhuoAa4+21Qy/yq7aBaQ63c2RockZzaf9HwmcT3D3fxLu62Gc+
Q3asjNQRLgDeeyVVwsZpIRKcnJSGrw4rtAultZyoSVTQokZu1FjsdPum3QdL7a3Y
i06qHgaTO/CP2+hN6uZIY8Ruku+420waeAUFT6ft434kcTIgbeLLXaxdiVJ8VU7p
vmgX7Q3VXihil/2idTDS2rYwQDcHYZnIuZ7zOpp2sH7E5rL7f6EF3DgMb4OBwkGl
sqJQkQqYDWwfQDTqd8RgOdBFaapFy5O/F/DH6Kx/jCwvgn1TnRaWodjPC8VEv50O
gsjx7N1IIlRQaX4MmSd9djlxE+GorLGXSlsSUmyXfaRIBAVe9eMzELK60mDJBX6R
mmavK6r+RazzXkP7Pi3MLEZhHKyuhZWMc6pkXJn1SaUblAbER+GgALDGy4/XcBWB
VXXB+C5FhJGZJXtdfz6fezNgk520O6lkwum+zlr3TBq+VxTJb4lmNQxLukgdaiHm
k8OdP/tlTO65YWnUprI6jg7ouaEjDyiTR/ejEpVeQL20SVuuD3PDmR65FUzn8cOI
klMluOZ0RgKtsdYfh2iTt1WQcY3QI2lyNnNa4nzlzsS6mLDej6iWrBT0XZiZoczA
biIvixujV9guXlTD7YPPdu8n6hMd8zUD/jr0eClpjrlprfHElnYN6LrcBJzvbxDk
rotRxwSxMqOqKdX2jk4VTzhVf8hmhRkjjeIaM+wmDOmLDaIj4LhjZOzTHJivJobi
wQ7x9dmVXl7UnAaZr2Oeb+qdO6Yc+VYcPP7nlXGyEW9kSyANwD7Wc80tuixrLCmU
JblGo4yoa1jneJEoPA1jBKbXqyOc+kbZJSY78mych02pAfQL81CPvm2kuBjIpl/Z
qO32Y1Qfao2Vteyrpj4LuAKiE/PupOdQoEbdpfc6MO5VzFS6itJ1wVBHepYoc1jl
JWh+jSLuprN1vY+Pbwy3K9Ud8kR1Jz7hKsRaIyHb8wORe41WzjyGZq+0cGpHetep
9v9bxFYR7vnyXdTMXzc72TBZh3i1vIQ4t26BU2VFN7ynyb6/CKjr5gv+TeiPzGqU
oIifmSJyPRXzhzxb9aji8FxZ6hPwVc74DtpP21EjAIUSImgClafqwZ01ILXsjDy5
ObA425aYyaAW9fmWyQnLBAAYclWvQ57D0qd3RvRFFhnX1JwlQGE9cUrRKgkb4MZu
1Y8xEzzKZSRVjCzFhsh4rw/lpj22OjLKBpNRdk4gdN+w9knlPRDbMzx4yI+doccV
vuKvxjbkrebsXSiXFKrclq+H/edrB8zeFUXqW/dySbkVYNXRoKfuAQ0Yqb6ower5
7H6vxcpLYSw1ZC/hLOj+yVD9SKDLFRRVeLRk1gI9SjE9ADGfIsjgHX/5W1caqTgB
Iv9bUX1D1upZrU1THViwIzf9ofJT7E+Sdk+thQBt+c4tNknAMaTNua0NP7k+T9p3
kUzUhLuxM4km1AAG/jW7qMWUddXz+F+SbxuxwBLmSYqkdW/h/6lEZU+qSI9YTe3q
iiq+qt7+oktYr4MBtRpnO0YlWmvHWs1vWkDVlmG42Iz7uI6OqNm41O8vADTQLM9H
9JlN/4DZMAIFiyt78pK0lD5PecLYxRsN0ss9PbVty47otS8vMETRKjjo6jP+VGQP
yopPCDkJ9aJw9vGak0yAWzdMfHASVSqS/2C8vQGYiIF4gO9Sxl1ePdAQH6BSB9hH
d61RaYzuWo0wajHY+aGPzUDbYhSj3SI9Yz+j23VUon7rds1+GuDlm7tpDeiWYwDB
TC8XhZKiIpAAeHN8Nx+qSgwG08pmbsafOwRbI+lOcbtyU1ClEupF736Hl9uI7Dvt
Qv+I8PahdsYqUGWyZ/G8i/TMxfUDyZUWUgx7Xyiza+KQpXr3Ri0NwoaY7lPilevk
QMwAU5xF4zMccEY+sEOzahhs18bYu16whMvxawNbzBWMrF+NKga9xuhXc/7mLboD
85gFcl8ORmPoAxyfnIJtUCfftLmaVtNBcvHBrg4Rb2BTe7NAy9SXznmmCINNWGSd
NjV6OYUW84VpGx+Ur+0m2PRNBRMG28/qNAF5w7dhIqTwN/ENyz2OxdzzhO6e3axV
3euOdAP8NdDHDWH98puxCFMHJp6gCbtaC9jl7+BtcaEa3unI1hxNPMJk7D91Mw6E
DsNwn1F0ZMiA6QMfX0FWDgzFXdXdNk2xPQJ5rfiQgtl3icqh5xqxh735inAXxvPR
aFgXBPTJ67j25KYycHCQq8+bd33YaB9BW/Ci6iWWWQWYnaBZ1dFyWD8cnmph8/Lt
wKBZSb065e8EskvhtO0ZQDkZ1UB6PZa9d27IPXPq7KEGyhkeohCzE5eM5/GZgZ/R
e6b0XTz8mlIn8Hwm1fxnd3JAB9zu4XJeSD9QJWM8XCVTpXfhdF3Ip/xtKQkfYP5Y
n04ELJZbhmdaYKE2ZRxx01HmEiMe+GDUSGufgH8XF6o6wQeB05WiO3kMSouqJcHU
AhgMw8prDbEMgB6DqP8P4lHtMwucc1CfHyA/Nepu0bCg2G6lMT0ky6AZhUUvTqkE
lcSrzkbn1/0Ab5Zqc3a9W+I9Y+nA1tOaydd/HPrJwEVRbzYEfo7KOkq3yG3FgFmt
XsVKrXAk70Onk26dzzE9sIYOx4woHwX4xgX4KgoanHBrcc7cQY5084lFPyBlMhOM
Vw0XodfK/wEP6a+cOCplTMqSPo7SpZmgLbAsA3sFeNcCHPVG/kWLgflAyFMvlccS
TZlOySaUTfeO+M5bsUlrnm9Catx78ph62+R6xprESO8lh5BBU7GXH6CL5CtlEAOm
fDBz4xmpWOsnes32gE8jYIk6mnTqCJTnTzIYPhTY9t/Zuln10Ak+GTndqEWdjv14
ylar7mwDE0HFC0n9/ujrCKQJWu8HjkhLhmI5+xxNvhgUXqOSK69eEXYBmIHLttkm
dAZphuY1DXyw9lj1V3mzT2qFN7/Ya8nrqcD3KGe/cquLh9YX7ZKRdBiXq6w/yoKt
e5HdC1Yytlo96akWQPB1EeQLSwth3VhB20EyAtSqCsGzQVzSegyINzfG+WXLvVn1
xti5zOHMlU6WlHtHgvkvyNYvcG1t2h4NAZn+S6YrBt9EqkwOBc0qdeze9HmhEmy3
YWqiuaqCNjdor8t9QL76v9aoIWjXDxen6n1dBz4Z8X/UqMf8T5wkzgKruJzZvf2X
rUJU0pEt3yYZQfKjRRS2JeRMJkofwAxSvXrkEKbaGO2ewAdEvhpFmGFctp/UZisw
tPu86W+PPccTtnqPzjRM/C8YwVkCRTsMmD08xjupd9S9ZrK2uSoCth33WPu85rzX
yoXQ0O00rxmkqRoqCsuhL819aZbERiaalZZ4EAfptGptWJDyMu9FmLW7eAxKoRVl
9vKb2+dGOB6tVzEzTrILitoduTLXki7JtpXUDd9F9930uP0FmnOQSUlD1CGXRu3e
3Ks1Eb7sLDz32BGtwuA6zl68lfVg0ibrs0LXNJsaOYkpMnhD+w3oZHx1/5aYj6J4
1/3K6bkORX6oDWzfHfsxInu7KLUlAYLJ9Z0JT9CTHTM2T7dz3PzGVP40oeweipal
ui0fguHtQqfYzxfNloXF+ZTSFByefiRZiTR8JzO1XBPNbTJN0xllDK9E8i95RL80
yWPAMDlGPYyjmfGsfZi76sHEIjD4q9WypL1XqSyFXMgfyb4KWXTVs1Z3FeAUMM2J
1NzybIV6mL2/VE4dQ1vtR6mJyDHmBn8VWC43rZxUz+RwdE4yfKgPwlCczzE0M4tg
oqBKf1t21S/y3pGw+YjTCT8PdacWCCXBnx6vjUqVao/PdFY/L7MkYwh/Cyw4evja
jiaeBPAY5LKOIfH+j0OWE8LQnO0t+LsmvOGk/A+Pedqs+gVUCMJ2GJYouNXdPyKk
w2oB8jKIIuZodHd3HDAd+ZOtziNRL1lrPQK808EM8DCX7LC8RzJ86As/INU1L9zZ
NXwqKK+PT8EPdfPWaviuluYlmMPdARZWENzUsfAFGYwuHEeAJuXsRJ8kigNM0OXN
EVFjR/ZJabEWJvvqoJEV3G1MTS8H5jbaYyekX6CQzjY5w3WohfPMXpdu1pbFu/CH
dZDZYUbz9HbGF7I3lzocF//fXlK5qM01/rFz7dlP0hd3v+QSuflN/349IrzYa6DB
PCGOjmy0+0s+l9GWyvWQjwXUmOMiHwbV1/46ajxTS9LZ/Vh6h3STF3/KHnTOoRUc
bp9rKpVduerVmgYMDborsGr4HfkQ7ahZzaspUkHYbeanEvRPfw9o+N18joQUVPuY
0H2BA2ZWpWTbAzMxoxI8f7M9ILhf6wcYj1TbF5shUFjqi1+ZIuPzgOddVmF2OkHT
NtDR3qsp9a6cEiCecNgKBuhJfqrKVTqDwoDA+0jsbNBxsoVyv89N9Vi/H/6fzH76
B8ImLOgkZUX6A+Yzctd3axVmfII5X9AhdYZryE5qa+tOJnby49MvJvtu0Kk8/grX
Rdr177F2F9Fps3n7lCzqbIEQ6FmTw+W0GAOF981onWVCN/DwO4GeAx9kt0z/XPq4
+0xPvrPyM0J6rsLZbwUWrQmcBq1hUSVQ5y+VAskJF5RSHfgdSHxLPmsl5R3IZYJ+
0xXX39DKP3/JYTSN0V+zLOuZHlcU7+Z2YARi5hNqOMcYrTWF4EfbbEgj7vimnYW3
sXey9CdkExOMYkgkFXT+TyONAlVgac+I7JELqCfHCTKvrz7iTvf/bAiNBCOjP2LO
end+g76RlFpVr1tixKXBRN76zrCZXTj+8LVwS34hk1yyx8wlU1h17LJ5xpM5ZOtB
f3C2R3hWD65EK/6Y2fg6paaJRzLdz2R2U68yEq3nvptva7KRd+8f0aO72tko/qEx
kPGhrjYXJkOi8djyNgK0Tguu0txGNsgoSy8V6nFgSbjf9umPr9cKhCJ2eGiDTFaX
9swJ+ZRQ4YQBRFR56lcOJT9FVN8K0+pcxNbQcSqmNSY4jEWyQ4WXq+DaoHOnt5t3
2MXG8LI+39XchYnWVCbDMFRuFCd44mD9MXCRxFicHK/+JaxQSJOIjqbvBXwtvp+A
v03eHp+Zpsihmya9JSbiE/Vwie+OG4SIzeuYa/PcaNJPNWE5vxnITp5S3tfLPBtT
iSYZhdY6iIb0u+ztWxTatVNajs7aVT/IWu+cDAapYJq4iIWPWmyPE+OH+e7H/rd9
XC3XujK+TkcD1IcUvMyCDn8xW+T7GKhUdEU1rxFu5hpPHmRUiaQM/kwY8BqbehBH
lIMqMkl+1TzJ+GUQE0+AmWJ6NQoy2CC8Cu3+0V0hflWrUWryfw2UaSAmXmYwnhtf
hFs5dm1N+V4RhGR0KS478sO+FmDRzROBTuZAAJ7Ct/y2yEuZTuHCjEqHxVgrnZc7
Dk6MKulInLeBloDKxL7z8q+LdH2QaxaT1IsxNe3TXOdxiiMX357zIP+VEG0EAvbc
UZffLqhC/fP7b4OkWPolx/N1K8DjytZ122QDB825Q8h9KpFq4VBewOmiVROu+cjD
WFpo0oEnUxc0Jx7Sd40P/csAcgOlK7qp7I/CN7ftb8bpQnSklcPrZLoFeLUxY+7M
hgwjKs4EZOPZMl/D3LV2+OsiO2cvK1mat1oIpC8ewAGj5A+265uml0JMHDT+h15Y
bPy4REhVGKPHrXpLHZZmHXsZKLUyEfLgN0waXRL95CjjoERZmVGRZdmoD2Fkcee0
ixJEcPRhw/yioYoIHICJ2makjxAMft4tIcJslx/tSNnaLs8hCCooJaNnuQmln7ZN
xkv0QDSWLfLL66jXMjlOzIsAUEGtnHdC+U7wfaRaVv51W6ZjPHwgbZlK5tIhhKDf
gxd9+AoS6/TNgsyee5WOdoQfbLm+rUmAYqC7dArZFhEDmkGeqMTXoCSmLVP9qOq+
ucyQoXcb8d0EUvKRuXQG1UnOsztzTzQxzdcrggRZm7VKUQmHL99ScmY0zCjAAjsx
Hka20oci5bWVM6U/0aZUi6YBFH7lSG5RivcIYzlA1+X7FI/SRcM1mfgKOwuZh/6f
Yy91vrpotcsQRblUpV/h587pd6fyeZg5hna3DO0/UL0EZrAnJEeUD8+3jI3accCF
QePxhtWf3RPhORuBknHIHaIZUic9Ov0Ks3TI7SRuWqNjJaqryouiGiFWrK6K5kfo
5xSV84PFV8nzZqpBaJkBo+rBFFa4+c1j3AVHoawT5oHYKWuRN+kmOnV2tsZ/GJHc
TeOc+dcmAlTkAmDSTwPm3nNxb9zoWBMKB4uPl4dCtSRTBGe4Nt7y1CATV4YaKpMA
CHFVFft9oo9gvpWyGxemQsddeg+JpNw1CuvjpjUW9zjr09jZpuC12iFtNC5Nc4p1
Kuwm7SO8ItB55EQT5gJQBqH+LnCZQnb7Xgnawi4x4wZBnYYiiPd+nUzmWPj6wAW+
2gH2PQtQkOutDdkROp9FHjzpUoxNzIuR6Ijsqf40/3FEmcdJrph+ilMnhOQSF5VP
svK6xyvCJwpCR9KkV8v2zRoRo1vsKEg33ghi13L+66m6dunj3+/vviplSoi0LD8D
pzCJnemtKhzezIS6oJ7VRpJwG0ajgW0lw9VNWB2CxEXGlkeHHugUVTK9v+AmWnQm
w9ejZ6IitPWf1vFWyOcqfuok+AGuvo7HbX32NKzj7B9oXpGiB9+ukJIW2xVY4zKM
R+HEYoPAa3QYn/3LNQT9780jwX47ya+pfs68Y6+z5gM4gnHaCpg3dlaBoOVkFYzl
xdZIHuORztXnt2y1sOLhb79DS+ftW59veu1a6edQobLwYwX1bm596GClgpd95DE6
sQc5BVgUQprnSWKGRn3avaNiEaxML1/Gn/KOnnABRg94/EqZSTZIeeNtQqdFuUdO
MK8UBKBQkFs/4WGDP0i5bNjiuysVUH66Oql6nK4hRHf3L+9lPcauauz7kxzAL0lL
4JIsEcsGxWfdP/1X6jBlKSMBGSv6EmcI/qia/FBGinWr2GyeJy+VNw/P2KRmqyTC
tbOZv6M+yy6KMOPLZAegRHDvS81CWKhWsgq8CFd04npSEGq7GYVKC2w/ZLUX/e1f
Emymp2UUCtSuKk7KqJiSYJLbAFO2RvjO/J0Eo6m2iqHSSmtHyVKnYq71sj4OsAmD
pDWkGz9SYULygxusCZQhPvXUfAu/EELUVa413k2Uwlwu2Uu9hSiw/QLxkK/+iqes
n7P4LYWokatDRJLDMQ2vz9+rXYSQ4CMI+wjMvekTVKotefiHGjZQsaWVVPeiaSAF
ZjJR09BiVhql9ssYe6CfpJE4k/qAFDo9yFNcl7Vlms8kdOL/IqhXw2LrN4nRceKZ
2Jxm0e5uvJGqe+HPidxJbeVHUGhHdreYug0lNJAgHXZeUAj579CuqivSzuJ3e+f9
TwvFMwJywmFAndaZe+kErpBLC6VqQCKTlsYHBvPwRfRQAv6TqqW105ENtHPPpAwU
zi+ptOQ68LiB22FmOmm2boCSe1+ttaImlKiQakOesQrDsqU42vMWNTyj4rRbqOvi
nEsuaySuTe1vi/y00CG0LtwBifBciGrFGNJKP71EJCxffo/XeRS3E7iMEhg5dSXa
n0NMR2/KYhjyHQtq30cc7okiA+AJ0mliyxQSLvNuhP/8qKwipUK7newODm4BsJx5
EyMmzeHhRH8H1ra+iAl8TqdNm/gM/grRLb1pDmOmas8hcjyL6P1aemeZudzzRN/C
8RM4qd9cifU59Z/G3SHPUihvl7pp9xox3bv6xUoHVFqGRUGuVADN3R3WMFcbn5Ak
kUtcSasBXAKxiO4axZIkQpBUadsMiXM9uPlDpAoo1H4hSOmPcnav6S3AdCjIcu3N
8xKPdqnBrhl9TOijYoNujq0GnR2AUZJyCMEhXu+YjJOXUdKFRhDqSl0/0h7vHQLX
KR/G68nAWzHfKJ5MmUPoYF6JIjLqbHz1+lElvlMdIERqCSIUOWpF+aCnMpYs9oOm
kmBFQxSippeaTAPJU8bE3Xu1mOfLr9ADaFi+56FiVVn5f7dH0gwSgtUX5vFt2jY5
IkaYnJjjzQdp45DYam2qEWR7kB45lp8pxK4XZQ338q1/sAh/+btY17qf7OUEM3PQ
sr3XmxxyWWLQ6F8sNynJiAY/1HbSd+yGMZDANBzIXHrCqrvJ1F/bn+pguG1Cq9dj
Hjv915jBUW6zpC31YnBZKMLnWe8nV8jnKYVaBmnUPWRYNIkrW4uuL72dFh2T0U5y
2q6CHZ33qwXNjLl/h3RiPFXLuiGqOilFX0OWJZXFC9l46vt0VZ8akb5gi5yv6T/q
FxWyo86YjnD9jVUpgSLCiORiq+zfzUwKdPzlHR8KucD8P4b3KnO6ampeyCngb4M2
yDA2gQDyf0kc8AWwYY6CmMqEVwEIYwDsY2BduT5gWKkQlFDW/y4JwZglkBqKUsyN
HVljpWpA/uF4CpNur9L1+xmZ44louxGY7WPBeOR0nHTci8iGFCNiAkrTl25BsA3c
m9ZVY8/y5FFgJYuOjVkQ4nkvH8vCTRiIC0NdBZcF3EWVfhpH/M+ofXoFG1guT5ZY
jhtqtUB2f6thEAXNrO4Iw8rGAEa4Hn4ncUNBD6x6yXoRw4HhR8SXcopBjywFk4QU
uiXoDiaWdP1Fig5mqbkaJlY6YKyTCWtahhHvWfydexxFIHQVA8souFbUzMccgnV1
hrpiNESsXXVIlHHxnKmeTIlGO1Hy6b0h6onaSmIBKWrCMvoMYEOCfPw+n9Q9rgJ/
tKYu0sZBC07KzhUi80lZmrT3Vm2u3/yZinXhCpd5oYYP/PCdLLePSReVygqozv8v
OmTSeJi3g9+Ibst10CgDjpfqc8GcEEGO617GvoXIzTlpKPDoASlUvFNJs4QlfGNq
BvR9vD3ZNsHm1HKOCxQgmnxEtVTcqjdlVqzUpXX6p1387AnaE8nMkAImV7zUvTtT
vBSgJqhgiuJ4cOumihdVU30i+g5E5/1utb46xv5XO5tAWIv48wf01NBzL+rEV6Wv
MOfjiWDDGV4Tn0pYX/+cTwqpXOJxnyNW7CvE13LOY0OlY9M7m5l5j2XantuUJkSa
jwVug3qf6ZGvD4ww+j+CNkY/NpkwmP+1/OFO93OJ40q/wwHoq/+X9TlUJzlkEaMR
BNT4Ibw9vLqttavFIxrRiCt09j4efEm9GAVpMcdSBbH4fegREIT2fs7jAKku6tr4
17dcDoEmjTsPCqGZvNaekqpplYzn+tg13eOjTw7w4oQs9Fxerosh3dhkOmjS17gL
WYjKXzvgn9NhXXlGrMtuAT7U0vxa6vvvJCW/WSJ1Oru9yjblxBRoud6Ce1ZL/LND
sDzmxC5oJubjU7OydfzEALs6dlR5iXy0ryg5UmtavFRMBUsOTNr3VpYq7l/j+8Hz
ok/YiGjL2ErLAqR/Fm4gz7s2hlgrd7aPELOFRMpYg3WQHNrCyNLky93S9wkFD3k/
KBs3mq1iLzLn2KxasudrLFleqyd0WatOQBZlsTreGQHnw5R1VfpQzp9xOgdXWDnx
56m7TFkRnCGhWN2LZ6ITxdJVTULzMJyqVj07RAYbcQS365SmP1dnQsKKrRTqtCv6
je86GN/gyjHTVjLBlzD0Rnd78uR+tu03lW5Hbna17O3Wbo8klFLbLSkZFQWv9W8S
WO9PwWoyvopsxghQq80sp0qKJp2KTMS0fPG0ecz1raDz3NFphtMzZn9HLStkhPLe
/85pCFNcusAWd7fOOW7561QjttkHCTNsRzEmXng6T1aSSqgnUoFSLxcJU5eXBiev
XN4cfIIF3PaK14gT9hxENZN9CXEZKDS6XtQ8u6JNA2VF2FUGSAnNxv/YVFzdl/QI
VrSwQ9tFNoFwwP6nqZQ5JNZtImTYcBUnCDbc1cMoy7a5AAYnHCISfvKsrfRtYkxk
OJiEDQ8oTcv3WCUlQMwrfqeAvcmxxwcKxEC1NUb+TCJbQkUzJQ6GjJTBB0WlkAau
BKioJKsMQ1wplKMZwV4ljiPDKkmnL2pAfy8c1ltj8kBwklTmzKOKr4dcZxMDhxN1
VTFK90sctZlJtvxa/XNdHvHYvnrz7/+3IJP5DEfxPJANoDti3UnTodjwKnJVr7BU
ZzKl9fANFZcuCeNRL1xix9mSbHGy0j9zIInYdvHcTppVHtTMJ5ma9JzmFUwXYRe1
clCIFOMSVw4JVnG3aDdrq11bbPCRiIaYSZn6FgsCO6WN+0RnIUPTVLKti+XWng+c
ZTPXlFCcK+DBWJ2RHkOtC71CxNRKu+L6e8nWNE17Yh7QQQVSUtGY/JNjNKeFQsvx
nj7c4fABSuID3BeVnS6AUFm3LHKwmwfTe6uIgEI0sSp/9byF1TvzoNqHZYCXe/eC
zlpmxztQDkFmIRE/Ib+YcYGs+aBsAMJE3eO7lff4al/Lmtr0ELEK/wwlyk9YLK06
Av03iD9E0jDeF13FhTTuZ6nu0rEDuAu2wOrNYxWV4hvLG24+4KkLtcMrbxRITO+0
WTTligXG2v+RFNP3ZrhKOcgCPwQMsy8tqZnysRRLxMk3w89MeUM85/up84jlI0Hu
JLPxvjZfBqi9AHbvd0520LYu6AnREA++OISkTuccpqwyTOYIxgP+t2D88JHOUSHl
A2fo2zT4eW18sJUIIZGZMUDVjWPQtmltov9LZr2EzinzwGAr8k5+1NgSwZ0q4WFY
kRJ3ck9jWQcRou1DzbOjqJ29NldUpBpWZtjOULWEUtwTrtDqVIe5t8a3M23fsWQf
bZmrB9zQKKWFZqKib2fgPE7BZDihio9B9siZiz9T/y1DURmTriKEmlMWIjrrkZz5
0hUpiGsiWy95bMsxLnBC5w7+4gkZOfIB+KMHc7yCKe56nSE9se2ffTISjoSQHFY+
IRIkScOBuRafy7M4gGlURIvM/FgKJqz/eS6heX430girSTKF/hPEUJrFkLSybr93
aAmZ5C7UEkkuPG0+FA+JqTMEnPBxnogvf/EWsDwwm3gBqZDsCCsB+0aCcgblIKsX
Mdhru04DWW1l0+WTcoP+F2MmgMgb4ceZzUaR8NYiSPzw+s0gi3JPTkTSpi+7cY9a
MOmuB0Zu0x2/boFVXYmwyCyqKfsaxZwizgFtEkvWpO3pflMmbG4dGu9zeAQfGFUC
6j65TM7Sr4bgHieOnfxi1VCFJQbBhmVFO/F2F6XF4vw1zn/NNshsbErmvf2M0/sf
kjHlV3OuhkqlVtwg9jdq7j9opZIwSKfMJPaVvL4FNQOspaDrqv3b9AgrlV7ZGNLF
JopMUU5kDvNRjFpbJv5A4XoFLjXyXeLGY3lO5RYLHbEAMS4ZVbnyMXXIQ6oz4o6D
8DW+Fr/iuYCZSq/GxfTG+8LQ/PNgom+iT26fP5eaf2jFnH/3pfvTnp/dgrQilmGf
syKtCuhfjLMSeyhr5r3Kp8CVr7o8pXxs65LqZJJ+ZRbvAs+WQc391AzTah+2PS6D
XmSK9/NbCrlVdbrb/WZamEwOljzrPJRuZHMiroHFrTAXDyEHpqsuVic1j56N8vTA
q5Y73U7azzSBN0xzw5Dme2IJ8zwQ5s7v3mY9PCo3Dr2T1lpYWZb5byE/ZQ1VG1is
XSiPCudWP1nnF6GBQ5S51U0t+pOeA/Xph6ZNyB7I/ddwQfnlwDCA2xNJ1ZUM1O5p
7F/y4EImDR3V0XQI3uaiaaVPm7hPRxRaTY4UtVdSXkt6tvKFbClj57+eLUtdnlPo
9IWkOPmw1YlQVkHtOcILwLvUl4dv55tbSKplxffqfQ0GmS2Q6zGX8Yk9dktAbZTr
zwXV/hFXUQxaZvOn8is05z8m++Gc+niOmmvLUlS37z+LR4z2cj0iyEWp7zkRgS+i
OIplvT1b73j51wj6wqhBF8gKWtW+eMdSgOB0geYfpE8VFJFf3D4iJpcPw9y5LH5s
HMmTF/PZXrxNOJDjddYkaMJ0xgOfOMkjMhSjt7KjJqDKKpjCj2Hj8+3MopFwqSo+
2XDpvQwAwAtqls+W0OORzIv6C5ZoFJuV49vfVyxyXe8Y5cnkQPwrU7FKDCMtGM28
wIv6yEABMfQK82urn7QNyG7d1hOXHEhO9C6HhVyqIqJ7OpIfEOeIlstO2bkjz16c
o46IGQoMwPi/EJ1kEEUz5ZAEwejVraAPgMzt3/MeEp+3A8o7e27YkC48T8FUeR1e
B9DAPpfifP9m365NEkcgJ17ElEVG1q0YueE4MXCSlZ8hdeKqxnqjo6DtvMBHowFE
yTTisJktLbdLTBGLxCCEdpkWUU933kS0kiyYE7JAPFnOhCcrESO0XPXd3dpiTrwF
WQiO5gmJAefUT69/W4YCj3w9YCHxqaMp7Vj39mHspgtZnyEffjoz1OrZMEwWYy5l
quFyVQpQJ+F+WOls4+S/py4oscRf/vu7YszbuxZ/7R0zacQTaDpyszbLQHbBNCHx
QRRIoG7k9hnxBmhZdI9sePMmscLkW04SfaxSekQtmoJNHdg5SsduP1duvBaOEytq
zNLlsJNzvM89Q4YnyTdZTjLDNeysCbEIEdrmfcHjsb3HidGb2ONkiL5uTEyFxxQt
AbaMd8uWYwrCIuRNwjneSzIzt+fo8zYVZKk9si/XK1xx/1ozX8LKWvFQKmRPCz+t
Wy9SWQjc/aj0U0Jvs64tpnR5ZpG/JyfyFzmDCBAZP4G2U251MXHv42SrT0iRzlxG
ZgUM4KFvmitVwexAH+yGYD2dgOTQR3RsPQE2yAv9KzMN8jfxo125pIFuYaADZMZZ
kWur3W6GFK6HLYAPZYPhqmBx/pe9A2TuERXEDbO/db4hwe2R02ZJksitRVJaFO0p
UuSj2pTXWXEeRjlJUzoZYlQKGjGXZPgfUZM8xp1433muy+o4uGfzuef+/6TWSea2
kfWCMUaG3++uvXp4aH4BVm4K0SGvMqoMy/GAjfPqoj1leTGd0ZcquowZUaEQdqwy
g08GKXG48mCPKqi6Urj7WRUTcQrqLe07bkmx4F7qOxPfwl3JN65sXJGVuCQB1Flc
6XGxgLuwGmsdqCM2fqVTWXfLe4OM2oBVVe2zPT61sEi9R8h4ep9WvlqKtBTAL/m4
LlgmZe5xOrN7Arq/sDOGVm1F0AI80NwMRdg1REfcbxqKBJw6VQV3oIFtlHmXyASa
orQMqE8QG4pjFJtgR9ps3CYTPeiPKOwWxf67Ffdo9/bzKuVPj9DqDNxObUyE4kLF
+ESHJAvYqY+vuUh0PyehbtMw+Cj8EhxbnBpxlzIBePGk2Wcw1lwut95vpir0goa/
4qvcnnRUTdtu6nkdZ/3xePB8OPaBXOdgUJboXW55M/oro62+b21VvSddflCI7FsX
qCAMzB6JFB6YWjkQgSVF1zvtVzD2iAXr9uq5FAeL+W5ogmXoxngQJ7OsiZK6NUXI
1MiFjyjaUVy6hMRLOM7KvBSPygI1YoG1Hzkhou7hGo7ZYpQnNObwzjVBQN1qcQZY
/JviTe875R+7pwrWn+jGN4UTJWHdXUYPyTVjDs8FB4lFiTK3AEqhPsdOl7ucVt58
KjkNfJiwy6zs4l1DE0wi/9885H0qvSu7bgg/ZHAvWCk53hwiJyud2RfIX5C+kEeU
0dOU1932sqlFRPYJPm6bykXMdKYCs/+vC6zpuioAD+5AsktNH6NXesazsR0IcL8P
8a9YfMt/JE6cwhex0WlaM6J7HFV3zux/cG26WaaUA8AeTV5+++q3tN1FFAabFKbk
C6GTIjMX9QSNG6JViEqZsBVuqMSZrWLnHL4UKjc+MahDjfTkcuiRCVryTeGPZiz9
KSCqVtEN0Kbj5dpyZ3KlMmZa3CmgyUr2EMvcFZz3hfTuNvqBSG02h2Zx/45sy2z6
7RB3g7a8KpwcC99qrUym3cCP9Wfw3Diqn1ZrqT0OYC9G6EOgJZforADmZ1HP5DR/
TbQwKZVHd2NAW4mLwQ3Zu/C5ZWzTHeTL961GGT+Pg8LMsNd1fe0vcMCbaAkm20wz
5T71FgTcxOw5TpZbBIHLsO5TtEM8RYQi3EgPBO6kv05KZiu09E2AFP/zmL0KVtPz
+qkA6w80w6mEkjAx5zF2dJGfmRswA8WFN+Q2TnSlolwhJxpFsUkuk825bdf/AIlD
bTr/V4ShiLDcAMJi8JesrPiNqwi6+OuVZHiDaRhkDoiCEhAEXrpQ91qbMgZiRhSt
go96hjaynig6HHpspWbNInAjpAJspUVnl59m5TsscRll1Dx4OfnOmhfHwM8p7vdg
kbh64WY30TCS5zjfLYZ8hskJpxf+tRQNorEEvwC9q2hQI0agho82lf8ibjYAUJO8
o1CnZ6bU/01O9Dmhws9aDGMS1VJKza2BfdEgrPSjEsaF6ve1dOLT5ZQ++B++JbTk
dGmtLGzTAKYsBGfSQQb6jmia9FrAn1CmDpL/NDfJcaNAuK+jugX7Q1rarQBuuFXW
rASO3o0l5ostBY+3/IU1Kl5Rmv8fGxuXjGVKBX8+mNGWUmOdn056UXI0kjN+p4cK
9Uwki7je3wjKbs+w8PmVBsSuphSlc0AtXf9tIEVrR+1FwjzljPfOHLMoO+gSFERc
KQl6IsbTC2j7N136yea3wPDIqlDwuNMKd1E35MCnubV8LvjqwdGs/ue3X7L4+pnD
wReTqvfoQctJeXQa6lkeifAvSLLMaZXLuq1uv7sykN28aZsMshdUljbDMOxPMV1p
tYjpcOf5FiKaWsrnUhR5VoGR8IiTISzBpBAnK6NMn6tcFi0ZyIw361vdsW0MbILS
I8Cy0ARRPOpuAnoD7vZ3IL/fJ8eKSF/IjFg6jgB2T4SGYpFCsnQggRtbpzMQ/D0U
bf7pINRM9Ru3TrK1LPXSt6hlahXRmV9HnMlwbGLVzxH5au7i3oFGNevAL/khsB9V
iGP81MgnXvdiy4286VsMrFNHUsg49gkfk5mF5IpKIvYMc2CbTgyr8G0yG4WHle6z
cWox0lFL4PGR2r1Jd2kRJF6e13DldrKaZrHrn8VRdd+0A8W4+/LysAmA1DqFZ4Vl
oulkyi/lA5Pa26Wqz2f3bmi1gHzHvcLDHfwYpduV8uWjQoJDry3l9S+jzyRTr3O7
82WreAtszIr/d33If7X/+LXxWf0j/LcHy709q4Y7v7YL0sbVitl70xwuqIHem16x
cq9EgK21ihGgbW5ZOEmSO1HexyCRzdaaX40jAIx9VjTwkvRo1iYsVBsFfnr1DR50
6a4TAykBQEAaXEnGEyc/kk3bqYAb7eY8bEJ6RuQy6JbAzjeelPWnTvLQrcvKVuv7
g65sPRLFXp4Cf0hHfSv/rxF0mt32SnlksizqEJNtjZe1SCxChekrsAuyeyU3MIqI
uo8kqmT/t+9Kf9eVCXD/X/OhlBnX+ILoezU7icYY++m+CMcRKdE6cjPkiwJ0GQ4o
aaMXSUAflfe+V8ShjNrLmQXF/UqNso+hxIAqHVx7jMqVKR7AvwE67MnaevAsMHnN
61ho3RZ3jTo04JuIrWKcbfk39wWBO5+ThQZVKLz/PtuTaB6h47W2G/SPcAZA5O00
9h2IL6rvq5MKdHFH9XKI+PG3Sf9qzaNJchjM/TwogxVrPh4WvxEYzkTSRz0EJZAv
hYHTaxWZ3+nZuutMOqhqXyTVI7oHnkLsyQCoxinzAmNbcjZzHVp/jpVfOx4Dz5tC
ZO9e2Q3KVI1VAk+XRFOwN9a0aqvBn0YyTyWv6FctQRHwD9YAh2AuKM/Q0coCLPVo
ifqi86iu10htJ8gmnSnjeKamYpE9ZGCn/yKn9QLbb6ItjE2+w8x8YV0jpAeF8NdW
nQTgaK81IvOFPwZ4ySOWDceGfcRt96ZhvzpvP4G5hBN23fzcSZVepftlZEVlyqzu
esjLTdroQGie9Kb4A4cnctL8t2R2BVtqKtONFW58GIwPJtxTVwiItJB/AnbXnHvb
5SeDO7Kl71mmPicEBVaq8Y8ezq6GxkwC9sw1hgc6fqsg867V14qzVfTc/OPXk00h
wRxmVQJKEfNiacZ4KCsmGbp+yLcfsmipt4KUYS99fw5gwe6jvugTJ8Ez+Nxw+JEL
9G+x3u+fYK1ODTRp/7u5mZvzzlaOlI+Y2zqbYq8EWP6XlagpH6EJ7KvA0ds4gs1H
rH+GvQ6ApTJ054qIU/7qd/a0lKog8sIZpulmAabWLah3/TxOMEpALZzs3BNXbFQa
ddNVp+KAMbPfK1AR2t8kzqAQ8c3WAN/Wv8PHxgpxicksh3NaNSPt4R6mjK6jCHra
MtnrxQi7Ym3mj1IXSkckgqMuVveyx0K9hfE1RJV8z9jJdNI6BmqX230N3vP+pW9E
EyzWfAz3Obnj0W1xDp4s80Wvx+xPodB8Yg9wseHJRiEScYxBZoxC4lFXmt3xloBF
7HpJE384rUTR8mNPEZHHzk4y5EjaFo3r9ys07i4XkE8yL2fkLErROJ41pt7OQ0Cd
n95xnYsAF/6+wa4dAqwiI6jQi78rwudUdZ1q+wnl+24NF8riC6i4KANbof9AY0Wg
YVVB4u86FiqLSuCAfhiwSuP2Tw6t2xhodUihBbx6GiiiYy0U9uIfhGO3yz3V3l8y
qSZtFGG4Z4JX4BzoTBZY6XW+Y1baNwzT8POPZHL35PI2UGGTmy16IeNX5UAqFDsp
Dm/1svoBpTjObZwJzQpb7mj6Mc31HyhArEKtbStea0qgbJFnGlsEACmiSJV4bfHh
cou6tINKajTlZJccoF1OavoMrJV8Q7B+UinInI7wj4Uv1MugJtqcYY0Mq1a7BUH6
pdtlAPtCd4jWhdYiqnOMcbqXjLeIlmXQTxTC0orsmiaSj/4wExpN7ooQcZ0mfC8r
1qPk4HxxOxM9WahOB0XY5K3tDwVKeEI7JH9fhbWFPIqllaoVXE/gthiUDJdjpetG
8Yije0jKBykuwe5CmcWWwQUTsemwqOXtOf6rVNOsvSxDP5F5JqwOAcI+f8OhwyBV
tLsQIGnfBFvextqwkUPEeJJd2sFTCwEKn2Sw9k5y+InJc7sOmCvXoGe3csG675O0
+b8ZQe7xM1a+Wjh9VHIS2QksWr4l/aewth8/ilF4O49xUZhszAy2fY5L+iOuEmPm
tkb9XZrZjWOAoiq2EYbq0Kg9zZ9w9nceaK/0aQ6+g0seF1B0S+Yj+zv1MCWMMP6z
7aee4MHY0IiJJYIkrAFkh2CFOjS7abRT5vFEL7F0Iw92NFx16x+UO7GvLvNzJlvg
u7mIQeVPx/H2xupBXgGbT69noMHrHzbddF1MtisxLts2p/PIEPmhG1ZOHkaK5YBi
nYZbwRXte5ZaSRdd19lVqbo1ZvLmNqmkNnnL6ULmnfso8z9NrmUoh2C0nXzCHZqW
Yvv/ish2CAC0COuxC0MyvliXH47V4f2dTuEKct7oLRPov+8Lg6M0Px/n3HWb6hmp
OBikN/IOrtuj1KiZtpKLfBuEcGZ37oauA5WoMTkJui8BIrMBJmc4D7ubLwF3zje1
HQf539wmBcw/NuAsgPXH0hxhW53hAyPXL1BjYGVxLwZNuNjFOqeycsdMrPJKbcd2
Ir8B22zcu0W53YF/ugRnN2Mm59HEpAXst22xswFTQ9mgEygQ82BbRTdbtNkaodiW
kRYxPcLZbFpW4lviILMhhkuLAiDRBh3g/aTGOU6v6syVPhdnLx4Gvcvsx5Gkp3Um
dTD+SZ2bign60iCh0JJawh+vLSJL4ckd4CV9/Qj5QXGK4jcyFyXc3dsg2Z5wf0L8
71cLAXhkW70KMu4F2rHxukeAzMcYAt7FoJNASN7IyVKbMbuBO2vYxdgljJxd73xv
oQ7Kg9po3KYXD1fWeHH7+flSNnkP9elZR8+VLTp7we2Nnx/S+JamtVzntEfWzIN5
0hk6fvtZlRrAEwTnNNCNJlCMk6ib/pxYf4H02s7l4Lu7MWcJ5LXyTdenJZDcsqlX
9y/ISb6xdc77sK/i0kuKDXq5K3pzZGqKLV+DWgxGbpt2h3tUhwztjJNtGmc0cv/f
VWl+hv5fqi+BR7bGS3pciZmB3mKT46t6gfcyhLmagdX8hRSA6la3nBTrq+P07iQA
K1GoTXaW3jC9H4B79T9wQiu83HKh/eDIt57oMWX+CcLFFlsPPMEWI1cOhhnasjK/
TU+7aHZXYdlg6DiKd4azy2mclxYS15p2tdPPiYCwb97uXdIkSAtpoUtXrY1YKVxH
s84WIHc2ZloxA8wvVAjxj9FGLmzX5GWJh64NNdQAJFn73/sNC2eF8bh9uhekd7LU
hhU/u8/YUFMua6n6WtcRNSfa73abV9i0jsSqgAxmPEaEVMMTMWYkFC1w8ZFbLkc3
q+P2oLACuYOn1Fu8vbIGZLS2D44AUjDVeIyUFYhlhF+wetJABynOnwa8MEfweTYX
P3XWTjuBJP9eArHhbFhd4lirSDcFKx8LGWDxRhgW2xKXxyzeqg5J9djDI/abQNIN
2j0+dzZC3y34LbG/SJSzsQB/y+ICg/cvbbio3iWYWLo6SnQTvRSJ0zKr07uV+4BS
fp7E/wjEeoVWca/Yv8jxYDpeiLvqpueFfqph5+J2NWLtLLDL/OfZKEKI/Z/OmS+H
5qxFl+16Ouz8w4e4wg+MF7nYMzc8gY2YOXyVTPVfONnaTd+xwgp3L8/EZTMDqu9K
itAlWSVTe1X+9Me06GrjQwUqLPRDylrnlamXgYmCeeytSxBD8Hpj+8tEv3meJlyv
mYDVsfBpoj7Pk/0SM9oZqMHNZuKOz/cslrUOT5WPCgryF8XL1xapIcIBBVid9A+o
Lu9a49l6sks+AmND1h6xg8xbrpvj7GaljKLU0O7ys2ZUdQsBWOD0hLO1LJjgUDv5
8wNu7KJkHZ7vPlZthSVsyLGKn+sH8zktTpyKSTCzx4czFn2VEAXns/h7oRdSwk+v
8VT/lvI9/pS059OSvYIthWN6R+h9u+1SQU1kxWMU0EbieOr3kmH2CV/06RY+dlxv
jnXi4J7+KZl4MMIRGHo4cegVmWIybK0tKR0ab0cPGjr6exv+b+bGUIvivaAkR2g3
NL2hU9PeHoNRmx3+LjxAFDOK5Z4WySoX87vsrJIhhbBwEKoBK3iDXJs0EkY2+eOe
gLfbSlxdV2ggPGthzzUL28YclbVhyf1pNRGqFDkblOcQJtPf9pkgeDNCkoUJOaOw
bDfNjPIQ+WGRsi8+hxgAKiisTHO3k1du/FKoorCVNUYc9pMDz8EG5j9CDVDu2Jw7
wg9wsY/wB/tzFNP6NVUWLH6iMwpSFIEr6SZqSdLy4rNCCDv30/jbcr/r2g0IDrpR
SpXhXjiRja4Pbz9P5DAylo+rkh78taKlSe+6t6BzwNxJMBA91ZZM6StubUDwA+c1
8+z4oB8GT+tHb2f/DNU9sakamUYXl98JqysTohbxz4kJzWsVLDUXsgfYiGSP6i+W
0FCRuYjwjNIZEIJvs3ahHi68FoWmCfwz8EB9RHgFHAp+Ac8xC6fRdXbMOj2ZJMUS
1Jwx1jdz1sbHrQqShBWqA9AM81L7LkpoEgzVgnFB6uCH3JDk18UVWn9Ar9uEDpsw
CtRDg2iqPLnSAwQoPaY8b9p/QpnZz5/F6A7QsTVLDjFCdgkV5qEiZgllU3EoteJg
0vgElVla8lG3sFLiTXLt7yj04LIfRmapEY4ZkF80xBkJ20dfUjAknW95gN39PjSe
aMjfN45b+MdJiWjVT7ndNwsmDU4cN+FtyEbWdeWqqTw9Nn9wHCCe8mH3Sr0QCq46
03TCOv69YzRdvK47tpX2z5g/fmFnHXWl58SxJIdaD3Hci5p+ysFgw4EgZ3V9t8gY
0sgLOT5ycDnk3DrARyXm2OkUAO7UKk3VZ4sqGosisyG1FTkcoXvlF6fAFE9TJzVm
ekn2WvV+O8uOODxV2YMCtfYwuGB6ZFCRnmO3WTXNAf2bTYFp8+u1kkmw+eXW7p5g
Vl0RzDOYP0QFLEPlGgiqZQetzHZbpzeXCWs8giGXDkFUVTb9X2rLEQE22LA8G3hs
RTSDXs0CBkfhM0tiafYPrbuNVTy5J/in8KuQDpavh8Xc5LXlh90xTIhszzTLAZSh
n2xiwhFYiyTgAcJU+ERvJ1axrnW3pqXpSS02Ci+bibDq/lFtsa8vye9+Yka9GAE5
Arc2RwYTnaHyQdwE9ybFOITsYozumruQ1nsK366piRHQoWUOQzJRR5JWFgVW6HkW
+Rt0o5kQpnaNONoG4vDXgjGmNsR20MqWlS4/kREQyHoLxHYwf9/Lq2r+q0SrlyAN
IlERYwoxorNdjdRz18QM67ggwYoyBj/YFr72lkEEayV72AOfoO5yqWMWMXaSfPk3
hbYCKh7Ov4zYVaFGZ/V9T7CwNLYGD27r1B/voIxXX0kyumrCOo5btiBFlwlnyIa/
D5G2Ln7yY5Xz1gym/apXbeylnaCSS/+gkFxQ4K1YkC3uFa7EoDeAztRKlCKgwncw
Ugag+Klp5xM3/jJAH4oyy+aBe5ppnraEHIyenD4bfUlClVlyKVUv4kQaEzFBW4E8
NLtQaJEP/LljYdaD9XfKl4gNIPsDJSuFvRw5TCoaYJu4dqWMGbzM6UIGhM78k3jE
ADIdjIAWir5/O9ZN8H+qKPbBIGvMZl1BuTcOw/yGw5+vOHUpGB2vARswJuTUPCYB
RIIFpG2qM1CNLbuXXEJwerhc/wE9Jm4uk+gUUCI3AbJNHxuzLWys7dCQiTfE92xi
ByVqwKc3XCdAy4/nbZJnjFBLNlcaJ4JXiitOjnDtxYNdPu+EvLM8YMhq/Dl9U+eD
eC9FEVWWuU/U0gCaYwBq2nU0Nsf2GYCK4xOoxxCKdmDew3IimGaih9Ayj9UVrTPo
yRbEgl7J+NCtUDK2fjo4MWxSQcRCT+VhhdaS/TRCd7zshnnV5w5KzFQaHvb0ndaP
VvSMvFLkWKg80EeqNuEUgMzIuMALuttW2GyeqolbsfzTTPlYPS2xOCw6jjWdryCR
nq+G2lfApmhZtb4qipisqByuCAP8QoAIF/mu1Dnr+tNgJWX+UeBxEptRhKBB/lYv
5hEyxkjkuZttdeVwnsDeODy+plgdiq8FOJDlgmn0EMr/hIqB8Muuve0OvotADBNT
Tz+N/DP20mfUWQ1QDw0AiqGIYYaW1aUQEcZ3DdguKyFx5Pn/rkJBfOCPZBd6NjyK
0vlfdVImHKTPxbM+CJncH5m3f3lJaJxPaMrSlyn+SUMWl9XNPnQiFDwuh/GqQHiA
qF4uaKhiTkFIbpWDaIM6AUz/8u6+Mm+Sr3ywyTo8YZHV9IpGzOO/gQCcZATIc4yl
qlIeYD7DVjbHp1+n9peNDw1FgZcjGSpWOcf7/gBVUWgo5Qb+XxN5u86bSiPhnYDo
Tzmg4QZtcRmd4y7fW2O/iKmz7vmwvWppv7pCXamwe+wzx3mL+Pa6+zKJOwMtv2Hk
dU2O2fSjgq7qYWI8A7jY2UGZdUW/z3vG2oZXrpGVUVg3dTU9zxAwlfOm4kR/Qd/3
j96yFL1W59kELVLkqmb+REg9sc69CtpsDv5WmaSOpetTG0XHGlqHk4+qO6enduNX
ARRc8kgxYUGL9wR0UZRorkOXBDu26bf+7FUg2kQjSxZ6/HyDBcgNR6ccASOIhntS
YN5hZd5or5cayeqeApXoRAYa/Jns/BkUj+n7l7MoITbB9228Xoz99Yyljj+sVRPK
1aTVgqk96vdfOu5+8geGk7+1wuYj7Kqlx9CBR1Hj/42MtxRXzmtJY5HAepUmplmq
uDeETilHZLHghI39gEep25StaAR+sh/KtuKdBZHN0ofR1AtUYQPWegrkPpaY9Fq9
Uhr7RlM2j+26AkBkTUvFi9S0e8CR5YDKN893tDJTggNSsLzHhC5/hqmjbmhsCl8v
6Lwqx3FMuufSjnP23wmxjK6PBp4oSZRLTyzxhENxiL6hRJVyLseMJF89N7TE0KQc
ji7fI14Qn1FX9rz8Op8hcniEY6e2vk0WHl4xjQSMtZP5fnqSlSuwbD0IVXQ6oB7j
uqqJ6sya/YXnO+qE0LDUH3Hi1hvg4rLFhmRhrCjyC9UVeTUU5Kmmyu933s3pnHuS
AHDAgFUyrWrABfEd4FrKc7I/tEIxuunggyfWQEPyaQXRDa0pTFG1jxglIiANUQbx
G7G5kG3hNpJT2QAsrUotuG2DbmMvNw0LrR6KZ6Z/JCaDFA5Vd8whvcjz79svJJno
Ou1K8y4Ry9kn0/jTcx7hZyJ/+RHqKrHkY4xmM4NdI9/DWauUaxFLl8loNiE/TaVb
FmmXiWFzjEXvS5NYvX2fgea1tPP3IOAW6RSMWU6mSffMrKg7kYa0X9wASdDnXLmc
DLjcof8zwnSB5iISyEtvIFc25WO3fTtHF3S77QNb0W+vzktX6Ek0W8VmGsNfnQeQ
/rWpgiXiqWwuG9KLt7mhZ7y7+JdRClHWYOJkTzYlniMQfCj46FFrnowpw+Ccmhfu
5Unx21kI/BC5Z9GdO6MHnmch4oVzcUxG8wjZbllVP4E1QNtyZD29Kv+klKpyWZmq
62ZtV3L7I8gkCQvhtACcCoipM8195xRgePbhWGPAfpc8Kv2O5plN5c54uomwJZ4W
l+t12TDUQZb/zNs8ZD/QFaWGh+3kxfGf0eqdzqyMUuAGVpKnY21iePmxjXehOLKb
byrmvXtzZRj/CbyGu0zZRx/sl+/+wjDXqZxsSKWFZqZghfeD7XPMCJ9wSdKgsjxk
TPuM/zTp8jJz8hyKLQvp5yso/yJ4bEcqwlMBaIjsexlTUpQVcMdNdIVqklCDqjeC
HYVg2+LslWmJxQQPcWvmTfSHXmdaA/VMsmINnF4/+J2C+I95g+KdLXd0YutK0ZZH
+kO1WNhgI2JuXXpN/Ko4li0HNKCakpWR7nLn1wzlaJGzaIZcvwm60IO2s/2hFSiZ
RGERo2LZPE8tVaGPgq5f++qUMlicwoIGLCgI1bXuYhY+wKDyvxhyFW1pjs6Rwai6
OCQzHDJWU0LSN5R8C6r5w6hXKuuk98yF8GtAQGhVtRcVRHfY2wMxVX4+QHsZRnvq
L8sXoJ+g05YxaQIk+xduuVlpGVPTZnnACnfW/vJUai+iIkrPMJvOp4UFyr6msYe7
iyO+krX4Oy7+JqLihEFWAPqTjLsMUrvYuQscG1yuKOSz6fWwJNYlVZpbswV2AnZj
XrlMNmeE873Q+s74ucoL7on8VCsqktUpAMf0ZfDNyqZnHjQAWNBZepwoZVzmCmev
5NyCdQvB2b9doVRTmPgl3cAnPB7j4WOPtho/TjZY5r91YF/qINem8i8fMy/cjIaA
NslB3GRSZUnYkab8mdu8A9O9TbA6CvSmbWBxyWdai5v1E6zYfNVBPQFoR72V1sHK
rnts1pdUbyLiB5S6U4o3w4JVVW8yO6OgpVS8unzdJmuwYpeEwgorHuNGqHi8+XN4
qPOB079fA1QynypTotFY/XgS6vZIgEWyAE4IoAmRIQcWaIrv0jIZ99MphBe8qgUt
lpjCU7veJ923dVct9iK/BGHT+sNomKm7x3ZyQH2u1sY4gQJXyE/tNXrHyBIFIsgo
319RO/ZbD72jWr6ymwvqZRYAK9hf6VhfE9qHUc4OWB0hPxjEinc+buKuw5kEUWNo
7ND2ah+ZwrJIW1mowvzrTOoiPRGA0o9SY8CowEAB+0gKcNXoiVFf20Wnl1/V8WlF
ftEtUyHAiaR1tF4PtPXV1p520iRXthdM9BnDUzVXMcfhd1+01W4S++nNldIxOCX7
genjldAdpgnsWSN27C8vKAQtq4UZrdATfPbThOA14B+XRs40kPqbi5MY4w5eyg1Q
SsSh9kbEkyfASDqdwy/pX2yZqnJ7x1U4c8nzVA73dqQuW1qnhog13xBkx+UBhSci
xNBiBjgypT4JrcJnOE76I9Tq1BErLs8865gpNwWiT0W45SkB6lYs5NZTEZta/zCO
FU8FDcns0YOHonR3TF/O5iQgvfHhIOLrLakJsRZHgRrZ3DPzzGweV62PpFACIR9O
SEQncUj+ZCx14I6ErJgg3qkajozAgzlMkI5qsF1t18yKAQjUiE9u4wzjETuYBjQf
Y41TLuF7nqB35OjtoHXyK0oaW5GoCJw8KnEz3KRFhenL1nCOO/QnFGEYWGhcm6/0
XFSRqiCqqG1v7/d9WKC4uwEy149VYXmtyRQoYi/j0UivZ0rubTE2Bo7rVZ0BF3X3
ZpchV+jvoupnrxphMkXZXzcExgL+enHmplCRSPq9sZtJ35eWRZP/gVeiSAS3Ph6B
f1Aqh64/UbX7GAa4poTbXPDYvbsu9hYPr+/R6f/tdvSr64RoSxG83QKzs+ltyVK1
fk+pqQEPUhhLyQ9PwFNqd0eKX4wJrL36LJcEl2Wi9LegIhtknmwx9yOJhFY0Ft3F
wD3TkjwWaSWmdeDmCKEEDQZ6lCFy0ndP3FpybhYCY9pC5sBAZZi66RAWBFGQD+Qc
ktPd4cjhFiq4JVMTFeM5APuP3oHKZnfc0O8KqLsetgnKD2pf0a0pzp0p8rxU1jGt
hqBN2dls9cCOBcRVuy+Hk5aw8mXgDGH4MppPCy3+4JM7QpLQTftwSOnAZ7Jvv9Nc
ppriOwoXQYgqFxUuVLKKeZcsHVqmk7sirsw7tkuOb6hUhk1zh8Hp9X7Urvn6L4Hs
CWOaqA3hX1mtWn+5+smsIHkOXmeCieczJbDAw2FUkWTc25LUhRJKJwUykKOLo6Hw
4C4icWrUVfIRGE9kfcEhYZkn25rTY6YCz0zhVA04HqjQPIslD2sQZSoYDNe0l0dt
PSwcPRz4U5+wek8fgIoSEkrZHK8sgmp85dZoPVR6h2QrqZoKH7if+tPMEPoutYlH
1EGgAt55zrzKwreidnIexE3sN+rnxWbGEtJJp8xYgzWKUEltF0a0BBGPiex63Pnp
DZ0ZvAcP4Xw1Z9bIsqFag2bP3QwlYiiIXit7hhjdUpmBs6JHTC/d+aZdE5dBp7Rq
TxDJN14xU/1A8k8D6+ddonDmoJ+cvR7RT5PPloetUaRUwnt0z0QzfUMvAZZ2kr1L
FlVjoZC8mZKSuSwLAE0v+4EhmMR5NvCUH3d6ys0qgKyUyHkiLVa2AF0vALy5fsTK
dCdxHjBnpkG673LOypnhl5u+0hGxNFYeMzwM9LuE5ZeE3PGDtrO5+A6iB/gumpeK
MAj+SlCg5EUVotOQo9snNP81DgfalnYTg0pPprcsFFOcEeQFOXRlMOhWX38aPnko
cbE8jA6wGtLlLXPECEaqCc/38T/nFYBIyGGb+mtz2eYN82dXWqrhjTsuEM8gvSta
8DYUOtgB+KhQpBvkjZ6KNvb5BEpalf4HN4XPbdkNSZasZF0bVUkzFsdHrf9+z4yT
AUwW605QTxqx3WkZKkLctJSkRz76FykGbK1l/JGLi+E/Hh0x6Oq9A2tj8k+3fU6T
cnF8p0LMBwKMw2WpuWKTkQblznbCbysslzBDPyJrqHi2Mo7VJdJqIY8a5Wlm8FSu
f4hTQhLjnHTR/IiSTttBP7aMz4+wvOg9Rjq6iRaKoBXcpaErkGY1bQOoZ4QwYkFs
zsdqG8yDlvyExeWrjgGYuoPmE3jxHPCEbiA4UJ9dJI3CmaFaHoxifJN/dmy6ikmb
gGlhnnaM/1Tdq/uc5Us6z2JtDCOoOBX0vaUmhTJrPeQ3/c2GdqGyKMF3zFomHI9r
ayqNAf00XnIVqEhD2SNqtmmxhzmBDwiAfzCkaOF3jKt4gN6o0PzaMyuQX9Q/7GEF
oP7iFMDs/4JK31SWyXDYf3EQInPv5JOJwN1xjlMbrRSc0Vt49S6acaKB3hukzlmk
SPBWB7ZInESFZaVFAvFrCgEW++oq2loiby+Y6cnya71+UaiqRsVqTiqUBFwBSZQ+
8slfWmfSygmz82/3WENiN/32cFq54ASA8Xu6CfV0YzOOSYIDWK6q0QQnGyHZD6nI
fpKf2v5u8a+X5w7grNXTap7HYY+UzrnIIYyBTqxT97afDDtrxInLwt8p5poDsfeE
TNwPRLdfX+OwGb4rliPrQn8u8i29aPjN0jtgNTC4xkMFKav4QMy/pFxCPGHrB/gq
nMY9Uwr24fHcs0Nt+ufj1bSL9cuIXNMJK9suCY7oJlNuwtrtvuV/rDy/Sa/uES/o
ha8oXTMgzo+DYQxetKm8U+45LhAd7TYNcOVWZjn9UyzF7VAJcHbOZjqjoCpX7Wo/
RsJyqhcYzG+VEXL6KNWLhkuRbKTX36uge0hwKVczF3mayaNg5cPRjJlz0HYx1jTU
TnkfPwaHJo28KWh6MvhqqipE3zP+HSGSZJmfSLlIQhR+oEKN/vRR7Uxfptfgxuzf
5O5J5Bu8sXl+hr0OUg1KVqaoKrRoI/4YZ9ELYe8RMdnm2/4z7nHs9ImlteYRETOB
a4cU+Dc+oq8waw9risx+u7wWrh/dL7zZlCm5XrdLY1t+0yPdsgeYmdTDOtGffv7R
h+STn6HLARAWAhR6gFcsqot9hRsHc5C7pk3FFUhNx0+o4GeUZKbG74eS0nLg+19l
HhPAkLO10YZsGlVRF/5F1W7vUkIeHRjLe3TfWcPWXXPI4CM5/uxYoTgvHGxl7plK
jxYpexYUmJXmycRHsFDIccNAiNBCLfr5nprPWjY4hQ9mhkk+Q3P3cjJKX+/8TyQ+
T4VnUPOVlOiWX3XFh1y9qmcvJozODHx2X0LrkRuecYISUTcnneGXU9v+kvgOD38m
bjHaz2n/RwEoD0AUPbBcMdUGZfnQXEmiVgJuDWkAvkZ93m9SLTcDgBgaHa6rG2FF
Ua0FtZjbCmCDLFJmbHFtbRnXSGPNmpwB1eA1K9U27V18togTNkyvyk+394Nb61Rj
ed6KaCIqxWL1ulMcnswkPnM/0WJik9rcU/AQr0cKNN+cy8fvTHpOqyMjuwhd58j0
jqGGLbKyrrvNLVOz2rFK+R3NZh5MoeRQ8TqNvTxovS87OHKk0ab3ov43PNhYuCQq
cES+s5fkE8HdDjocAfepeuo4OXoU99b+URev6OThJVN83UY7aVvYKsy5fV/oB0Ze
c29YozmRPtsn9t8Y/9Yyqzl0yPo6Tcd7xCnL9tYbNTFPffbPw8XJagF3rfZiIctZ
LlpTZlEc1Ogczly9SGt6jfDiOJ8KDOYi+P2xLp0dO/XKtMi+roQUJ8S/2PpysxXi
rLi3g1/WIYXh/DT809lITK0MYSkId1R38WJeyuNAdCZLCO2CyYDo42/kVpGwZi+R
BqlqtkDcRUsr8uSHoV51LRG2weMn9JGv0Rf/+IZT1cc1aISowizeAbzVf89dcPfv
6h2OpEp+Jmpqn7Un7m74HpGiUW4itEOF6zDbEW9WQhjN0hFqLLYbWPJmvra0GZwe
E4elc08TlGTLrH7giS2CFMxqa2uQEiu3aqBN4m3Ubyb6Cg0xbyE56Pj3nZOW9+gE
/E1k0oPNZFRfwBU6AoCUewT1cj5Oom9rFO1DwJmRc1+hOpTU8p2YXnYnAtI3wC8S
4/mtVu+qrFe8W7uE0FEpu08CXXaef7IDPUbppfEJl961yhoBtgNKtK4Dg81mJqqz
TOTWJi16I0wFEuqmQ4LMDMi+2RuXF9tLyOh6EI+SxEuE/LO95qRK9pKutGHMm5ow
AQ/XW2BidTWkRTj4KyIAG2fnejJr5pK46+3Xa6uYhhq4jkcz30SfpZFnr3skEfLQ
wio9Y1kdC9LK4BLprKuQ4fh5/ruSc6dpIFT5++SY1d5uYe/eyZN2EA5oFUK3Fzra
usx56EzG/gkU4a89NuB6a3aFULs7egJxe7JR+DT5qonF6IAmekhnbEwOARlNDePw
e2xme1D88BPGiCbS4QEXkFO6yGt/R0/d3XuJSl5nOClFWKc8eCixaGk/UuUbDiYd
T4yTx6ayIPZiBaZU6hGY2EbYQjn7kmiJg9gVBWeRLVfaPwb9cdkvMWroERnjiR9t
YYVWuu0BnpKJlW4G5w3n+JjuJuNApsZ72yYYl8KEbbUvu2x6efYpDvl/8qv1ijOD
m2BTyvEAmavbEwoRklYxkqGUrC82MTAjsYe8dZwaa9Ft2CTtPflFa2d78QMRwvnT
5glHJqfFw3niQbkrn15q6wjTSW02ttlbuOB7k7TyaGsx7I743kMKfAHneB1DUDFf
XcSmmnsTHskkHaPlyc3eRaeU0W+TZzHXF9eiGHSnhMHdVeiGw2cKqCd8sePrSVkP
wGvmI1LClXn0zl0AQadZmZMGS61Fx9GH/dwOPFoFu+XatjjoqUW7KTMY6EyzYfb/
KzOWbpLXxS+Qdg5KU4Vc7CXuEPFwn8RNK7JV0jdyd+6QPWWEhXEHu5ZsxgS1wLln
oN1edJVY8Xrht0K7Q9BTM66ZWoR0xm+Oly31gIwsiAqSXjySCLN1yntDdHOkvLx9
3qEDytv4hZkVaRwGil/SuxB4AJpRANiM3jA+izuOqqtuUYzwQKoe11zB0yTQqwyj
kp6HWu64yXbBTEqyIz5Mh1DyvXRWEC5ep59AsLPw/UVhRB/8NIjdU6YAMfxQF0QT
5uFSO4b/YCREX7PHwlqSXeI1PZ4wdehqitskUDYjSQlZDqBe1ueWqxPSAaTyrpyN
XXnnUxS3IWxu6dD0Mh7h9RcnB5biLyTO7dsS1e1NRC8lTKxnRVMVnVM8oHXxxKMU
aIlePtDX+7Mfu63VQpVD71NjpyqjqGgpjIWa/7tW/nFRW8vKKkxxBw67FKB/koP4
9C3oheQF3oyX7pbzhat9srhX7IbFIP8PicZwQxfQjqiWP5DGQp1fNq3fJ2e9KELk
Uo3tSQSNj08cDBvB0O3d7KVLShEryiCnlANS6JsD7C7bR8Kc+KBcEJ9s0HqJv/tM
3HyWxZRZp384mg20NJ/HpG3NYI7XMmQuaYEqkPtI+9EveZOiyaNM/+NXiwe1uing
WXhbHO3XePi0/OLEPuLaDzLVXJn3hv/5ZhmOo6xGpkKyw7nUXxTZQT6LKe3bOqfR
4D/6g8AAtdQRvaMnfaU9EkIaLU3KulOv93bU767fFBjBjMy5x96s4VVXRIWHJwJ9
QpZa9siyY+9h29v0sp5r3Ikj+n4X8ReXwX2JY6p5AEc80PHc+ztApI2fXmFWpe4l
lWlxJn4SwpOcPnNvOX+bXuwPDA3vv8yyON1LUhnw9NL1v0pyrtu4JqwAzSQuWnDE
mbuQAxpaSFJ41+xNLsd2PdhGeEvV2GyrD6Ptd18AFZf/Q4Ti5OUtBYTdgzc+ehYU
KqE0x4xttCYRBJeFM/E9Ab00bvU6dttjjd4ViOqUxTBDM8WBQjuo2TyKQtNMsmYj
hro/NHz89/mCchEckWS+QUe55ic0dkZbjj+w/6IMLK2AUZxRutjX6+nIhotJFDys
R4JAqD/VCBaz+H4A05fitwsmmG82iRw18ZvPtiEm+LY1Jd5HsjjgxHZgrLb07614
dVvSc3cu00rtBaA+BGXLY6rJZ9v7ZuktHvd5H5uZedf9KFG49FjpEIobDbSUca3F
TMhKw7huUtsrefUTvIEYnZn1+NQKk3/wFtHs7q0QXfu19OdDm/PL2/xQTnoMhsp5
W3T0GJQ2HoZ9k8gyrkkE2YBaxCqYdDx4hfouNMNNnthVnNaM8jy3cnZewauIBf+F
kl1ruIAqnwdU0NYJdQYSYKj85Ii/wHiFHKmbEEnjGVUraprjKlZKCfhfkb89dZRJ
ieE/mdkocqMfQLrfFUrRqnU0aDdkPVTnAXIc1L10+GtBQry7cLo+qntkRAm4LpII
bHDCICe3q7DZTj3dNBzfo3iiC1/uGbhRHCwq9BtFO+XrKIDc5h1oqX/HkVfWtvxx
JRp6Vs83BCtgXL596xjbLTrmVIqII5Z8qZ47viHkQIFlbUHcn3OuN8f38gyif5TT
xy04nxcVp/fsEiPyJosZaQdk4gcmUYUzLJVSDWRHYEvsSd9BqWuHmoH1C7j5wo6d
xU2xhsKud1rU2ioCgwLi/wbnM1maxrZbi9wYn7A465k85sZxL8TwoSTjDEU3ML2p
ANN7GWiv0YKNfwY+8XSLfqzweegvda+B13l62DZ8YanA0RsujuL3yORdjpkB/AO6
+IrE5ywJ3GKIBpoisobsE7ffyancawxM98mKpLcMdinhzxumJiWeFVFEbrtIRsuj
8VW1tk/5Ui8EhRRr9+K4inT8yfngdYXL5xWzwdSGO6tCQCmzd6FCN/LyKcyMLS8B
68HllwzHYAnELCa33mQLwO3MCf/PGUZQly+7TkseYefE8roUBnHvGHoRI7/w4blC
FzqV7y6dt0XGyfCvjEuVwDN1FTcMohFeP0BPerZa5S4a7PCHDq0HIl1QUtTAVPqT
ntylk8ZpEByzla7mzLdxqdN8Z4FZYt8+uQhv5T59FajtuL6qG2Wk83mu+LVPaIhs
9lE74VMsRNcGeQiCCi35caVMCroI8co5Gk/z0BSbhnq67cGfDl2V+JJq+t7lU0lI
YjJtbthv+aig6dFS6ojhmI8PrIipB41BXyj9Uf8GE2mtNIKtOMinC/bYCvLDOkSm
N3ctKrZwNf3U59TgjA0NxFs2RvPee1Cxh41LCOFd3bpJZDdYuyJONVNKAvKYZneB
PVSHb79fCZ4i+izJvsJHCSM/MYYDrg7TCNRvplH2T9+vwjgxGJJBSrcIdIym7CzG
+tTZOmJ/tNNxf9QJc3suKXO02y/2Jmu617pJZ89ZI69F80Ys1w0J6bGkFexSwme1
F02/Gxp2buoI1PJp+8Mubtb0auUgfvCB9n9a/Kc27jw0h+r1lUms0sxgcwNdXOiB
oJihP9zjAUVNN/LjjQVbS67TSxduZk8VRKYp4L4xq4icy5KBo0Ph/ivWlfPKTF4S
oejV6B8Hp2SDlYTmVUYZe+Gxho1azn2HMAQwLt0DeXNMwTzPXybZ9p4mdFbB3Wlj
UQ/S/5UB416LgJHnEfRcxmIz4Hkkl1S4kI26ysT4afipmPJrpD2dpBip7c+CFWGJ
YRw/IA0Q4yF+kQcg0BL9q9XqXgSqDO2He6mAgG2l2H1jUrMFte3FSMDAxfXO+J9T
NKB9l7wo04b8Japa3eYt99ioerP4+QvtWJh/6psIqjm5OkEUAP7t9ibAu/RQg2Po
TsJDTl0F0K9MtHBr2P8fWx/2a0KcYT223Y78cZMUI/uAEPZ6LS/kUtfAAApJU2NP
yQ563r3JGtn7rsDFthVJbgaJ8V80fsgO/+PM08Wj9zXt4ZfdsEsFi8oOGodAGLtG
XwXzGU9orz5N8fxdHFuvmuQH9i3B/RROVCxpeWUU4qKydr9yvi019ItQnPF1tsOv
FT3N5nQsQZEJcpNBoJHE6EGINRkoAqIFBXGjSUA/KdzwnyivCu6JJpKgmiIh1CEl
oU7C4RlXbCc20/Vs5HVLpvWpPaJHy+wO8G8NHp696dP4wcm2oP3pQPM3R5+TOfmr
RSykskgh5g1RHGv9s28jkkmdxg4aQ5vAUTyM9QdwWhNGWnILYTIxrREOSgy8iFtR
n1QKZJK3s0T8g+oLTnnZYxQncW1Af4yqNAZHisBwZEbc3Kbl8GN6Zeb+dmHBuR53
8qdxEd6YbeGxlZ2jYO2mgU01iAr5nSj3oVor4ANmAF2QmVOWlkSpnyTUTP8gPlRI
titXTRVB0w6K+J11HZhjRNBwbG/DLvZecgk58l8TLaavxjnihsxtFRV5kmYp+1JN
Np0J1bbkS7acMwxvp9pyKuaRbqouzKQKkHF1tA4kEiB8tOq5H3xZXBG8M52tLiyH
yfNqODgUU9rU9Fh/owI9EUoqW3BbdPjJRyXhALvPQYNPq60ZHhUou8sGBRCF8Nj8
n2XYMWel8sQ0J50Kofinqry/SZM/2u0c9bClha+MXCQQiKIj+s6vz18TnmRNFAKK
LTufzCHhx4x/Mha1JNFHuzwx8wk1HC0aCooY6GODc4D3+LJXQ76WdHHEPYpvK8rn
uDQHqZ6xJzN1vT6DnxQZijDPG9JAHcZvgBltHxHyRZwO6OCeqMnM24wyP9311XVd
OA/YUg1AzXkgsINphNarr5vAaP5nXGUlgwsmEStGjDSX0k0xps8ukE2+K79t8/Ic
UkEa/dUhFIU1IxoUD5FLZD8Etz6Z+4ZpgjRlTY4FgdaLKTRc1iLf+XNnJPyg+o1l
s3WFYK/lKhiedIH4Ko+521FrJI2t2yDdq0Ezzm2YlMOgzPq4hz+bS6IS5CGcsSpT
CtLhU3znYlu5YnWG5U1DMJ/mcQ3cp4uXqUYBzz6zqDHqzuoTgLkIwiCIXmryZtdl
9LwhHCaobPpZMwTu4xMw3dfLrrVTH42zlV0b2Lixs09nRWz7M26eVz/kK30ZkMcg
C/f/uplGbjfwf8b5N1h0fWxQqTYExZeOuu9oa7HfEsSIy6G8psi7Ozto4pnJ2OgQ
SFVlxvvNdio6sEPlF9uO8p4LcfVObe+XBaS8+WcM0XlfXLgkRjez6li9vmKZSfmz
KJaxv8lb49zvs2Kj+jNAd4RwJXeuBP0r1XjAlEMKTlk8oNE9jS1PCePavjeDLxeb
JQ76061BK1yhDAMYmPoldYqHzWOpJaE096MOlcKdfoPYDviYUpjq3dX3RTK87mQt
dysCoubrnmuCBIjJLltdlVtEnx0XwB5gtokbc1RzEiF6maao4QJ1k4u9zxZZtm84
91hQTgUE9awKboqSR5uGwyMKVJZxmL9aSenvYKFhjzqzeeb5ERNPcSuzGAzF/UkY
91tKxhPlPxY/w5TojlVy0OboVL/Jl1LQH7ehN0fw1f24CQpsls/df+faJYVs+N4m
Cj8nzAsQniqoCxcwgm/aFFPuRagugbxp3aaY3XMYGvnfvMSsbyOw58JOwaPp3meq
Y7btlJrQ6GxDI1DhTnrJtUkPY0ZLkBiCsXObiNU8aYTkSPUG9kzOqSwrg9VCm5D9
j84HVkYdrYO19KhYbNgqDvGz740IkEOEuyG4vISf+wzbOcp+aTIzCYtH7GE5g817
+3UIKcEPobJxRAZVSAYbkVb1xXVr0u0iOXQ/u4MUUeI6qbFUbYYGqMRjNvVgMt6t
BDYhf3muXWH4b287R9wcGizTdgMHf8zedeFyFBySKsnd96226+eYDo50TyFbXXJq
ucJyeO1TK6CG6ab1LeKr9WgUdnpVpqWPAgQJ1xRj099IYNLD3zYubmyc6Pm6UsdY
gE3AZ6XNBcrbT7ZQBhq+R8K+V1N+ceVql7bcCJCUxqSMzlWfY5ultXcosTCyPZ17
T8xQ0s5vTSb6KzhrQcz27qVHyDlszNURTlIctXRj/Fd1YDhsvjMuME3uovghIjJL
EzVCmZ4yeM/NU4So//qhdQvGqmK02HxcEh2PjQDfOfsZ+UTWUsEg9ehowEpwwIew
FN1eblTmxfMcmtpwYa9qKNHc3lnt9vuOZ6/4PJhmlAMbFQGOfV68IHY2nyLJWvRf
QNQbiKcvkJDtxz1QlMwE4hGxJC2YH6b07xmKH7AbQMdih8NsyagqNDz8akG7/o+z
TAptoGCpwujn3iMp+scRhgd0LhXkNzy/oOdHlVODkbF2UBCjhHDWYGN27W/mEv+5
esq3YlNew+jhDjRnNUm3F0lVDHODwxM2HHHTUqWkan61tBbuo4McDdFbmgEXFtW/
/X5XMCzAXuaY1UxCONZztc1XVNHLHmyjwBlQy6B081iBsl4X+1ibuPgi5Qy08ctf
bzqHRDh7cgtLlj3jFmnncBzR1nk8O3LgzLHjS2JUsUzEBI04WW9AASEQDH1/wjqf
Hmr44QXDRTF+DovQrXVq7zJmeFttK6D8FAgUcZ0vU1Pgp1+/ia+2X8n/zsfKbbd4
sUBcbLfqJUoki9iY37iiSv+W+o57EEBycTpmAB8jT5A0hwqW18KTnv93QteIKhjE
BD981xBg2s1h00mnfO3YFU7DKY5enIix3W4XvR7pvs50GG+rBIacbis5ZG9KNcYf
9fGbuy1Vgu4YpkLHGHXAZ2N7b8M06hGZr3Vd+XHRGJ3u+/8jis7IR6mNlyQKQmfd
DUKQ50h6R73iqdfrKtXcFTULKPxrqEyg4/lO/96z15GH1mfs8D7BWhXvs45+Sa2s
ZmVgI5mEk2zPFR8IjfUFxoFE9T2043i+vj5VqYlRJUVhXTTcixdh6hjtzDF7HXUO
VqFwCOUiu/+m2LEiMtgjxdKEd/mBX3gPqjj1RoGQ/pOd17WTC6sHo7/ARkjm0ZOg
lwxPV9IYrELBbubiG1ZPEJzC/UK5LV2yTXW5pLcIwBqmsvMsXDWmSubiPpW4dCZm
h83AY/rQlk75lNgIAGzKidm3WFMfi6cNjAU4u3pwopdoNv0CVbnuqtWeflhNFUNX
jgAJIpS3ipCL30rSAJQNRrZs+1k1BphR1MeqZpBg/yZDhE+PSP5YWfuJVfW/zNWb
gpIt+mdz9RysG7X+i80bsu/q+GJsm9uQPSKWzfoI7F5M1bfolhnolBumUUJTLfve
R0rPDUI5LaGR+otjCj/A1uwbhASKPILHZPiLVy9woBi6R+QO3gG4ZHTWIIFi8zYV
uQqkKqblE4k44PbEAVFOboTNsRqhibRcKg3YrHwyj3WskTspmVVB1vWimmFJ929o
IuT73sWcubfUpW5srLAHuG9Y44G8TomEsW52QVvlhCrdGplPU2CkKHyTq0IIJTmM
yZzYgqem6APmEK3yZtOZCsjwpQ5NNXrb+7SrAjDr7Ew3ihMzQ4zuTDNwY0wRuEQL
n7npRVR6EgCQryZReMGHaZWHbXtcWCrwB+1s2bxfG4Upn6B8fXnkIBFUiG3BraYT
k0146dN4G8l5SB+V4sVw16dwn2HL2sHBEIU9pisKmKuKGE1vYxhfLNzfWCQLncZ+
pvJ2ExpnzQadrJ0GiUJzmTLyQEho6gUzqArEUKcWiTb4BPdE3kzxVbA2UVpWz0MV
yJGR2vja5wArUBr4JomXzkkCGLG7S2gxlFZBcPnwvcRcylvVYQ2DtuuLHz7b7J8+
v/vvIa4lSUonAWrQ1RkYGPHpADBV7znd4wXQbOOoF5dJMpmYWoqHStZh9NsqJuhr
BYuizMP3QSxs9Dg6cyCUwFjMPkBokgj+dB5YDw5JURfdu5D2dibauGAwd3LOOk4f
1V4YAEEsb6lNbBnIWZEgJhaGgwK4OGFrRYNuQXUFhexG7r7WdwKDIsAhrHP1CcGH
d4k66X0KTeAcE/RvQ9/TirdK2pRcQsNzZj3sW58JGnQu1Ae5JiO3tjCNwMw1VYAm
uo2nVyH89f95F+2u/gk5YTN/d0R+hPjhnWMYiHTCPDsIpUu3ABaBNvtdn8ZAu+9k
rYVaaDhVZCYsMs2lgb0XgvWblCGS8+ztEVHSlhsaXqQoztbiTvN3KybAOrJ3pqSy
cBDtOSRPwq2Sbm0bsDdJ/TzNDUMnzMTejDlNa7hc1Xepg1oRva6THzeXFjYU3s4F
glG8o40J4XexbruW1pmNvdEQOsuFA6BJpUj4M8wBypBoVI6f+KvcvHI8cLmgTL52
Kbs8VmlT4E7GHJpSYU2bbZbSIpuuhl4xQbVWZUsX16yW3Qdv/vV2bwGCoawUGGum
itNUQR9yq8BlGPq0qsdNR2VzH7+YFpnEdhaxuZKQ/rIfx64mua9o/DXISQK/caNo
cLsrIiiCAtf4KAOdVHvOhX2cqNXnhDDKb/tRimJqrTRYeXCY+ksgEH1mGCevtilE
To/e72AOCvAWZABcymPeBWrZwsc0pqtQ4t7xX6tllCNyQCyZUnkZDqy1zWklifkb
msCYS2Ypb7grFw1H4BtfHbnSEfASbpN1L9K7rpqg9o08NNm3pljy1AKPA4YnSgWh
+LXMLy1KUro+SA/wa3UqnyznphmVeuH8IXsWwDQ1hzvNXfc0PxYXy6XUyVMtZXKw
qNXyakSrAr3C5AXLPlaDAxHoURYsKTqopjyLGWApIuTzpfNlPmmesSTn3LBCl0td
d6L4CcvYSCrLfgAbnvkj+Al8q6RhsbNUkXAoTD/B8WF4ohqPyNNYJ/AZg68LB4uT
soVxyhXSQr12LIE/VKtNq5pIa/A39hrwkzvnwfOnjQhYepwCpcHIlI/7CQGA6bSL
CZDoa8r2Y2vsXUJW0hSjLAPhHzGq2hYT09/ZyKuf9/wv4Bm3GorS+TTmlVA97WVi
FXpgDyFPYGzG0khVKW0YKJIeudEWSjHeOx9m1T8ni8uOCpWIb+18AjhP/VQHStgu
VTDgDmlPDDy6kFhk2ZOTiibRHS95LMhYDJuv1eau+v64yGodPy3VOO0ng3CvyFJi
sPFdRSJ9crlk5HhQ5+BHIuL+OPUFmeyd3vM8HJ6NjSFyW9tVUqSj2eR98XovOSHI
IVY5OnEbVXW8snHk1Eq7OC0V5yhFCLAk735UWogOdOdguIWKmGkRFs4Q5r4XZYYE
3INaNwSVlEwZlJZ+sCMQTM36neRWc44iz5ud5F+8JkKBDRkxy+fj91Ys3f0rAC/J
By8dB6zBbKA5ZFNndk9QlBxyVF8qpLAJ1CP12IdGwylB3wA/yTl+xqw8at4Ng2Ou
kXNypB+2p4dSNI9S8y+tcueQKsH27Eck8+IR76ZmmKRYsg5Dg5k5mHY2yUX6yR8Y
8gR+4GJUoRmeH5rSNDgNY3m96ZA5LtAP83jPP0pv4zRI8fMJ1lk0uwvomvqvrjlJ
E0tNuRRgVRInRx18xTe6WQ/67Nfus7juhzFtQ7noXlm/4q/YflBUI7qoRQGzsqwK
V00NkD2cwIL+mdJGg0k70jVtsLWPrYu5CIhxf3VFQcDAptbqb6Lc+HXgSgHZDLka
1KZ47EcUznlk3nVt/jvBxXGCrNtrSLjkOxSlYxA98UibszGl9BM82ddhrR+57EJZ
048otb6d2cedIEQSAYUUJ1Wow1883a5jb4akiwnjInMMp6CVB7UZRRfmIl6hQoTO
ZZqk9zSQVmyHSa+6pf/oj9AwSOjPdj1QfgK/q40422OiPDjtAIwtWZOYW98kcZKO
ED2F+OHPdMl8mvT5wLDe97Jj3fs/fDt2NIcP9w4tf52wcfj2U54RSkll5cxtIB7q
Qz26eUN6+7pajXc+Cw0wW+M7l9JQjhTM58PRE8RxAdyQkIZC47NCknUfX7SMUVpj
P2F4cHeGAtDjtxq28oR5IqjlW9HbuH1hq0w6+Noere+dtGjWHIh9SXT2P3y4x9wT
nhbeCZw2agHtzYTr8u9lhSy3qhN/Ukh6FEYdCGTLdz/kwkskiUMSb2xZiu4yKHaz
7b4LhvKZeNo0VpG8CPyJDfaJDNMb23L15wkJbZ7CMwlaFagXFiSdoN288J8AcirM
OMpfSacBuC914+wGyKIWedYcUEahpc/DKPg4MDXnNqEcsBDgSbQLTJRac99G4c8Y
Pd1GxPSAMhsvon3UuKNO/IcO35a+ed19sHGCNgj9+0upGQn7vmTPXo/kNPq2FyEP
RHsQuFbgOnMUke9J9MQ1yFJ8k4rvtYgQzNvQ6rdDf6jOiw61KlOogh2gdQdnYS9a
PSssQnuU9yRTdb41Aszp+EKcEjRE2RVkC8+DggBEbqtx1Emj47JbUZ5Jvjg5d8nm
z11PGLFUeDET6emopjMY3MsITSdWBb+pXLKurjof4/CKQ8bdEHjNTxVglDMPN7W8
tJhS12EP8usnFsn9ElzUfA8JNYkUhPk7byxJiF0PH0hWYO62B5Ayo4z5JCMtdpyN
btKboiSylgvPOCrR7bFVv/oS/qsodHJ5i1Im9p3/BV3LtOZt3sGfDejccFaPOXFf
w8FxT+6BZXxn6GPAZbiEQ5GYiBJ+BeudcuTkVkuWM30Rx/knDwPB5wSZcsCKdtFr
prDz1f1drJ+Yoy3jfDajrhWpjLishsehrg4q8af74uwiVy5/zFXOU4SLKV5dYNCm
7BaKIyGGCL3DhQfCcWA8kLjOuHb7PX9zL+2Ic52Iju17vtBv4JZhijRzFDyn8KAr
Uo68YmW92MSx/RYh0LgNThmiUP/mxJqxB71LdbdWJzw4yZUHPAHA58j2WTnYifHv
ceMDEMpQIakLqy14IrMhekcSPEiMI0uEeDySFcxZ1AGclQ1IT3DJXo06yQpb/7R0
jmWPRzQMaxWgzvaVOw24OwSgWGhbe0s3C0VAr9njLw0oLbQONBRIN5zxk3gLVbcZ
GTmOpvh5OgoSaP0QNW+kPVeQbiv6KgbV6xg1Q3Bn7rLlEYhWTvXMqdzqBOx7k5bC
rxNX07hpc1lpQY+f6yGnvkGcU4LO+8JCXiCSf/lM6rKe+jWDuPUd5otRmufo2tkk
KHcLbOQwZ4LvwQxT5FULbph4KyAyyfu04Rbp6L0tF9dB4IpGUY15WUUNXxENZzTf
EeeAHnnjour9R3nApHXkQpm/OfnLzKKTR+iszOaurqAIIs8b2m/In0qtN9lFr+Yu
XrbAu8gSMz3uHiWAI5XyXFmsoh43doXmaF6QR/QyT1YgQ6jmdS/ilYUP3opfcUyE
0/clGJsITyN0NsmUXsf6NkqIFrjN5kU88yiB1eG4t5wFVuj+QSGPjOMK86eafulE
u6C6TafePKhRV9rBEB4uC4FfNQBZyrGomRvSSY47OpO3q7dO5bk29AU+Y1OiaIKp
ZrgsY1+rhOmhnRzXh7cyXsGhz6T4fWCXh6tFTfGAus/JmXcsNnEAxfMbwIT4BPJx
/wnekobR6vmTy0YRnDkuEzsCfpvv4dT3ibdCsAIu3mpMEuTyIKIMcX9DphZ6t955
2M0XYriT0iT0ViGgt2QKTGg/RSOEIIem4TL5gAGxE3IP5Fgae+BYS6rMCZ7VzyKN
g0Qic4f/X2dBNzz7xcTY8vricedDbKbSdw9giOmgV6GrhU7WrxJLmvDyg4YjC8Mr
HpWM+3IN/V0pfF3ek0wpfG3xNRPem+N+uU6EVzL3HSEoGpRHpCMIL8BYGaIoa4Gq
BJSw9/O2AUDizUw3QFzYL1HEUGJctmVS55kfjOMUhs/4590DCPcysLgTVTBP0dFM
V2Ze69g4t0yLpXPMX+1fCfHydDWoZjhZQ6sIbbEtIb7nW1V1OC9kIkOs+nNF9L9I
E9WCtv/I2x8Glev/AuH4NWerNDz+ORUsIorYgoAcExVevFKhiDzt3N4crlCkTN1p
ipxby2igezrtrq7+M4DKjTsXbe11EIHeiWK/EwjIQpSJSvjs4MtkmwLHX3YRq439
DQ1unmU+buXx7PjAdfnU+KrAAcAPAv0URco9Ju8Pa5IEiVakhm2u88bZadRAD5di
1j/LiUicOLFdFTvCQZvvNuRxq7YjsjIseMhswEy3Uh9Kiacs7vkf1L8UoVcSNafK
SYIT3sP0TyrojAqHPrIsB0bljSSzxh4uv4lvihYsFrYE3PgQR8Jl6WDx3Lt+l3d8
4MHpfGMvdekSghsWRRQWp64Wi8vZ1S6ZabPAyftPHhD711AHLU26LaspQlCZUX8B
9wKIv3L2sD7Vskx7ZNVR3syrcESPAolnFBzqoTCSPO7oLk7p7Q7Rk+Fn5/IJgW9E
0fUMHGGs+cFG2/WH/JxS1CMnEeosuEG9K12uZuca/DzHyfR1DPDNJc9XDxnJd69W
oEZB7LoRBmjPIA7L+WJSO35AkV5fOPEDeol7Zk/QOOgHnqPF2IVwLYQffmkucasU
CXhsoOUzX8N10+VCSNVGmGzDmFq3aad+RgE+fAcbvWAw/FguHxEclr2GjCjYgIcj
ww1KlBNRYo4eVXUi3ZRCXgLj/mWmOLnHO/pU7fI+pSCpore71BCUnbQlSEVemQeh
lokv4Kf08IJvatj5sGfVtUw4wtfWZn15bQPCAQjJfZ3VfcsxgGzuMsT8yJRujeUf
YA3E9qENUU5kvLjixgT9UE9FPbiZjy4n28OgCd6CZ63FNQd8fSZpor3+kHLIXjci
Ik6O7H0lAtC3+/8BFfaw0l53QxKMykK98xPXXHqm33qoivsSLw9No5HkV/TzfIXn
+N2mUxV7W6dAHH3ziuX+CxMqUTNXGulWQIOBkkUGnmxGa4TG6W+u6awBdoaO18Xm
TUXB47Bieivqc8fHesKq9ek/9dOUT/ZHF4pFnIDme0r1CROcud5iT4pzmERDZs2s
SewwSPg2zcZv5+MTShfjJVYINrxQNf5Lu82ar5e2/xQBYuDG26+zJlPcBtNWxFXB
J3jlg41hx+p6Vu3PZA69ydW1ESra3eIChG7x22/1nE9h2inRBoD798zdScJ5I0vu
VFhdgmrjfYGPSRLh62wrUhoXFGUUbor68g0OyGUz9LCt1xhfyGRCAq/QzSRxR+dD
S4LTW9sQNrJGlBkZ3AEda7wlD78hvATB2SQLgtm8veCsprbvkHM//K0cRZtKlN4Z
7ZhcqEZ05Z9Xtpgddm5B+KwNtunqU3hL45yRbMm15SkR9vMj2QM8mVxL7YvOgDUc
KNCI5bF16auCUcHuOoL3ihoiXMB54zycji4dOab5PJ9ysutZSN6tKzHVTpGgaGN1
pXpbofvvK2tur05SYPpRaIBYZRPchomidtEA8nLRu0gmRrWbihtJWZoF++SMWnlk
qBfBxo8p2zwC4SSg07iqxefNwwFHJ6YCHbS58rRMRextyRoD2r7ezkRyzNNPa/6T
SZ62ctzFuvMwAY1dU6NEop1D9tIz6F6VhPwCBzFQeOS+z/aXixzNqA/3d6900DXS
EZF+ap9ofULynKVUlH1BMkgZwgOXZrYCIn98FM/e1PmpQc2SNzBY4/KhABN+6D0h
VAit+ZxmnbgDFkq95sZzU5W23WXydgWpxOi1VwMv62QZDAEoO9AP5fuQZjafPpAH
VkSoQacD3Pj1BQFXkZTHqFq5rXJmabKQOOfiJqLUdhkX3nKEHHfH1CZZ/Ikbmlf0
A+tIpOCQhp66akSarnXpoeGhzREPCnzFuLUyMG+kKg/fUH756OiMAu10uKTjtdCL
STdnX65n7D07JD1Xl/zSGTUUEUSngiTOs0o7UAU933uhOWOF56Jo5ZVPsc6S23o+
XnyRTbMA81dwaJgrXPPA+1lwH7mANe3NKPz4AjOgeP4wmXQxsgxz5YDn1w6y/pVY
a3j8hAyy+PDgcEE8fnYoblwDCoSxvUVWilUWkswJcfOpd8zWAdjvB2VxJwcl9QEW
GOBsrzm0Y/CTjr2PUdyAmcHFZfXLKFf040WcbGvqgPlVAkbwgoJbaiUfD+9/+huQ
CSe7FIKQ9dTT29N6HwMpYW9oqFkpKPwbALMogZ+PrGEQInq2bD+eSWbhjFlxatDp
HGsEg4L826nLSJpH40BV/wJA7MHqggCxOSaKgljYkstjGKYPm9E31WgFDxcVVHE6
bgXtByZeB0jqSeUNTdfpTGya0qZxcptRaVFHaDiFOYIQ9eywWOK+w9o88aG+A3S8
n8n4KM1rm1x+hT2r3EaHg9hGrFG61kZ4Pk6DbGIN2/EdilcSAIQV867bnjw7SO3J
X+RJMsXiVTfYeet4q4dhmDZ9uGWSNH4DtdurkvxLvwoQf1H4BxFV3qcHSlZwfqUk
rfwxJPCgXvLJPhok2NHBaMRfMlYVildbY4ZRH/a6lG6UhdGvjhQhE9wKsyqKwO/6
jQUTb4L5VlA3y69mPgVjs7HkrZz5AN/LM/lUkipdZGtYu2c3oibU3z+pN4pgQ+jJ
rAITx90sKv+h/Zy+KX9bbTbgSHinhTBx9RkTrk4NwKWDivh9mDW5ht09XzneWFLm
j6c3UUzOmCXRVQpSNxOtsfcB+3SALpuuWzjCyIlShW3YD3S75JrhEdBS9Ea12uU0
mh3FoKJjg9YUU66zPD2/pC5RkEd47AY8qIxdmskxOoRjuRUPeMWWgz+eDJEvJRJ4
o2gbK6izCtOSGJ6fIToZu20FCP+XbEhWaRGWOTG7cxzyciUEvPiXYfjPZ08OUXL2
od0gcTJVE89AetEtsp3aDwpIalzyKFWjBwl0fz1fYO1sMgEsG+up05cANJf9EcLH
Ud/+X7FQiXxZQrBRuUJQ6svrgSgenU2jci51SfbmHGPg6TfjdwlaRhFrV6pFAyDK
6u8Ljv+G8SHgI2PcJuVPeHJE9Pfw2zYTSq2mGLDQR7mkCwmGDy4tGf7P6M43H2Pi
DP45FlhZpJ/J58cr4+Ipz8HK6IdURWU6LqeVDFRvZjoItooBnNnMBWIlxgRnD7lI
rvfMvqOvwGEr1CWJ7WHNnwuwl2ll2T/FKMz6MutxifB6isQDx78vJQOBQp6FtizS
S6gnkkhjzoOWaD/Ox3BGkGdaYeikWa4IMcHLTXPMTmvPkriQekEZ2vuofzYUAed0
Zo5H5OWecB+lk6ziBJuZz029D0CeRTKvjYggR2yN0vD2yr0Gb0X1Q8Ko3N303xfH
Dvi9mKMlGNWljcZuGSBo9oOmgNLfR5775OIAmmSEyyZodQ1ppJWId0+WUc42AhJl
wlcFrVNnhuip7v3/Y/0O+a8Oflbjmms9Ux3J/svwtUlmL4yGwGskDp2RlnBQ7+AJ
125GC2dcebJa4aw90sAbYb2+kUwgsxE5eePSmSkufFxRXywfFBPezD94iA/EwjFy
mR6UHrtNoEEHvQiPYO1kRZHrgJhZ0+kVJh56D1p8vkqZG2HDv/z/+n42vHEMw1kd
V803OQwwUZWuwUbZeyjs0NOCLObQc0juZdbknzlA+4malcIvzJ4mAUdOTUOMA5g2
2wTLEXCrFEnIOILrZKah5YovOvkFGZbYKIWWgc7uOOx3r7DZbC62BZAnzv+hczCX
32V5S3BKKho9BHEYLZ9nioXoSO3waRtp8fDylssOyRd47U7pYklgDvMRWj1Ln7JM
igMFaIpncLuiKyxsXvArCfi60lksuBn4dmUrljNiOfHcSnMV8gglwzXhVKlZJ/IS
wg8YrZuqXXxNqgefvIfmBVSci5vb2GuoDpwmBiMN4loEfJfqbnJ9VIrTQ70mCfEG
1/Xk9h29doOTRklPNu6wX6lnuWEX40WkE5zQd9R/KNCiwjgO7Lg35ED/7ruzSn9+
gB6eDuWsr4aDc17Ng+9PJeu+rutnOhJzUPJNN2t5ASAfJ14uo0pD3hevZHssRPyn
/RwLX0t4S5NYWGjAz6DKI9YNn4Af0fVeFk3WQ/uB+Y2NE/ccQnlenLzJQqngUH37
vqbCzkYVnkl7Gvo7lya+9A5Y+MphcjNFJuNBeVNna5CN3cz8LbNZAhzol7BNBC48
an+zYK7Yo/qdm3aQascycLgyadt1Yj9cSaYMKKlRhZFOP6nRzqBJeASkG6isH/bZ
LJ30E4Kp783roxvjRz2OrEBdy4t/zquYFMsdrwJu/2b2SP30YGxx26IB2CRWmSht
qSniQGRThvRLJCH3MJX3mB0wgKULkuXVuXmV1DaMtjC3A2oVtU01+ucbNIdd0GkW
tJP0GdTvLkSO3CEgHPlJ5BX+hXypGqY62PTUPPMNTA0ckbis+wULdtTJ1INYliq0
X0gpUeMj3+ph56R+PJ2eZ9NTz2tKErs58KIYAOAfVweaVeoGIiV23VpowIyhgEJI
EFMR0glJavnrKmphN+miFs3V7YA/eCCvHoj/7+kWNbUhgTjg72aQ1jW9fXoqRxNb
IlOsbfHRQKWdqqK8KHH1sPs7AxMZULbiY2cklZ8Q4vJaWIERFdgS7356LCmmdS5d
b6vP7c3EQu7NNziiNLPaLrehbrG7B/IqPC4YThI1PJOMO5nIEbXm0qwdzPSlkJaB
q4Ah8nyRRyk5KGyBnBdoRB5fak/QBsvp+ie8gvHg10c7WQX8Q9uLyRtlK54PLtQL
t8Oiu714oxRSnb3ib+QWwuCDdoeqAsgRnjDR1kASplKu14dQKuHCQ4zqCBpf85X7
K0Z90NbYMXOifomXBG5lo5iEeEVd2ZHew84moNF4ltHln0x+s2ng71CCY8Zs5U8K
+jdTa41Q1c7E5mFcT4v89jmHJ3is91rVWxHMzXW/woqEyOfTt/I9aEWLaG7yUA/B
O5DWcgc9N31JRQ3YW0XiT5QTVdQkd7Yq9bQSc9qbggFCI8dhFHiJZaqipb5LvAPt
g4EA+nxHRl3FEMW6kHg21Sdj42w9NfMyEOHMPyxcXAltkxpxGYYXA59VeWvhIpHf
/h04oS89dd/60Bn0GOsemeK9mIAx/W4n+nz+W5KkZQK1qQRkmrvEJlthJ03USjDd
GWO1ZU15HmRDOmMJToV8gVXOTTTvcwUI/piFrDz6ONE5h6UKyRUJ5wqmV+IdxFCd
emKX+AUZydUGRZMIXRuqxkP4azQu73t/vhgJXQd4ZLhInrU9pvY282Ned3Z4toBr
ogMpgMbw8yW2nQu9yM+fXVRVfEhI4IxbEo76QhtuBaaeJo08j/lWoDAViJm21Pjz
I0a4Zt922FbwUfn0aC2MXG3EnkI9c904ow9FNY0X6jivWtszhhDTkEMVwTbqyg3c
G3m8u2iVcbOhlpXAUcuKM/j6W+kgvyWTgGKCiqfdjTxcYt+A8DyNcQyah92p8XId
l/v/1LOEoKLWzJwbhosmUXZSOFfdLli73WmtNfzZvuM7lQxKhu21miJx63ki5YqY
jTy44gF4TR3EokcZ73J/atpKYl8GijHWiEF9FFJfGPOAXxaXHGzbd/AFoLR8V7+1
33xsA3Nx05GykLkSfLu+Dd3gio5Uuy0uRylPViYyYvpbICwd4SI5ja8UPeFz/+pd
5Ba3EVxZ+Eqt5jUAAr4tANpZr1ZYlCI9Gxpv5pzsvarnJgwOua+5G07Nu7/J4QCP
/URwv7Ss60bDY2xpWqEHvR/6bnAioMD6m3wstzhmY+BAH6saEpvbDHFFg/N14xK0
BZ6JDgSBYWQKwthcQ/xuxQIuRGRjaxHgqWcMEfp1ph8hAaY1OYAfAaCQxwyhE2tJ
Dh8yPDn6JbQck6ThS5DKnetHPNL8jVwC1b/ILGmEoaEL96tVWUF3dRkzoAi7rs35
HhiiMGahLxFUvdDHCWxM1aFttrafbXwD8a6G3UfuEp9HQqILRRHHDe6cYY+OCngJ
NaROTaIZgoyowTFAwOjTuc2VXJlOCF1Tc0liMkEZViZ3p9WhiHLRBLqNJdsXBn4H
kJFj8u5hjOxBIXa+NhhSKGex411mEd9XK9pnSzgTk1Py5mEm/oLzMGqExgrGT4Xs
mFEtJbC4ZJZVrGr1SAqBV/nCfPqqPzL9Eh6SLxib5WfRJbrQpSNi1T0/e3hKX2OR
9JrSn3ZHg3qsdMb4Iz6eXMFZsMKIdfyNnSgV5JFtL52u4EXZ3SBJBsW8mISeKnjD
4QyQteo+DGHM+gZYjfyr8xdV3kRYgJwUzz0qADY+5fATauEe0gOh7U3UivxqSZ7C
7t3OOI9//DoIo4P6+CZq0Ma3DpasCbpV0UATi7bPrRj+m9LIVou1Fi7JHwth6y3T
La94IzyLEylGHtUwH1zGnEpFFjXKo5BcYZe4d+diuRg7+hrgV5ds3N4dN8XxrAA+
Eb/yq2mWLr6uMzkwNwJoZv6ytpYR6Zx9zKda0pG74rueaTQocO6aMXC6Y7nlG1/P
ZijWMT59b8jRapnqo8axW0WUSWiqkdMjz0gLbQTR7OjkRbAoTmaS0rxMbxNQ8Lta
kXy4YMlmrp2tI+hOWf3QMCc0zOG4R38els4JNI0CX2RBMUNrKnP71Q4kLKzbAuyt
HdRtDLIxhuzxEEj9s5hpm2yFRrr1g9oorUY3WFOX2WuD9GcS4m6SuKSJTWKjn0qv
7mEAv7hvEXBb28tpC9xJxliC+tyhVSFjFgPD2L5Ll6BFjY3mTvyygAI6P48Javgh
YCwp51dAsqr80aeuR3P7dBteGsrt5N54uc2uAiikQPv6B3ZUIp/Mx5MwmeNuMGgQ
NBJLLY/EKe9DYaWWgJmlk4FbiQ+rcpxJzs96jnNYOw25jCSLj4D2JMH07vxswdWa
sjCiBH/nWcrSGktKDAg8RYX1+wUgHT8li32aB8xIKysqJyb1BxkUNBulNIJPWUtt
nEB9nbLlD0N8L7bG8Wc/zkH0zQD3lO3X6NGaN3MqXh4byJgdezE4bMzTMouiAvkF
23UMYNa1PH/any/NOJkA5dKfvmd0KNsfftAwqul19dB3xJFTvFkcLmO3FSe96FE3
pG4KIrGCtsId9o6KUddxiTML1s0+fim+tjMweIqKEuNsZN+QSs+j2ACvmOJ2DoNa
qH+eQceF3qxeSSaZalECxsyp1+cNBQetEnHBfq4S7cVgtk0xHTU/Ft6bayBdPOf1
qZkC1ygdVVax31hsbYS1DnGc12/AYyN2qYJ46HGDyvODvlyXh2RAKbpISiZlFVLb
y6j6ZQdifrgnzxOOs4QphgMEsFYSWQZx1iZYHNdQFuixSSfeNsp0uO1qBj9j1pS7
hj8WSdcUuH/XxQ9KhfrgFm+qH7YD8kO0557w5W8/3aag+0ocSk3oD3B2XRtm+7qX
iJBQHn4Eg78iL84FhEqQk3u83E1cCL0ZUSEPKNAsTQWXdcxFgV4GS0bC1+WMaOV4
bU4OgPEVVbJD7rw/oSnE6nLxwr6rYXRzHsGDENaih/xLJf5qwtw+ZfVU4N890ec6
U+7Ec5i3/mPkClT6eObmLl1g50n7RbBqm+nUkRVIlK9xTgEzqruGtncXNxDg5wn2
4P0GUAXArYhJaf/CxGb5+a1wVp6O1aJXvgCDnBdCmK5ACBIVmM1WWdfYH5H0KXiN
+fJ+3fANwFLCc6Zutd3bKPkMWHpO+hS/b631rRgWeKQEXoDtvAxSwYdu4FfViHYk
FWi2Xss4zSIjCM1zdZeXl5e9OT+qVQ5aVY6PWTZ3zAZ3eb9WrFa6Tl48cNHU5ZVc
DJdYyit5VDyQmsbn3JgEdLr+rpvVGM2gLoxFH01aAG8QveAiTDxtJEHRVk1HVsWP
LxeOe/JfYYDxIhH5AIJpLEwSOXezoUYdfbyFLoYuDgtbT0/NMNBhKlLsxtgBxFMU
F7MgZEZQk1PMW8JcXLpbPT8Mo4IVyTBcJPXk4MmQtPT+gg2TIhWwk+LBj6qA8B1x
PqeoDJV1Gr3KzPF5w1QJyAszmvS6WHkE8TI5r+w24CY7jMNb/TEUPwi/HtViSera
vb8aONF4cexP6ubypS69w2QUo25YLOLXAev+q3kWtPxwmJ2Ej0ENGkEmkm+Nlxf+
uULIWaY4e7PcNRLemtDOOSB6Xgygni962Ie5a4dcoN8gBs4R6UwUixkACrjD+sKk
T278WmOoWMBeJlXE2tauev8q8/2UuggZq81p7y66PBKEcivcaDPnUNShL0rqaTLX
BAik5qnL2tCI/VMkTAF8uxDcjJLtS0rNFNcbY9jV5nfSGAH+sXhjpRKJl4L7/gWH
o+HKnz5ABdFszupbZqSti2XtMxTS436lsH43EeLAZtCw4xfGVA7P5NETpzKbryHP
45R4GB9d4+4KRfnyMGr6f2HQ8baBqP7ZqPS82O/y0bta9zTus6Bq/2g/Ud+c34kV
WXUMziId8IzdCQsZOA7ATjc++J1WsghW7/r/n74nlwNdebffSed7CZhnmrrf+myH
AnViKXc/UlanH+/6LULQ1gBqHkEYEHbIciRcdfJXj+NNY/2cgkY9SQQvQ7RUqKBT
BtgKugUyasPsAuWRBJ0z/PSTZP1ONdprJo2eyg7lgpLeBTOdhBA6hG41avPPGF6f
qwq3dx1dEps+jUUymJFGHJ7LsBcC2waa7q5H9Vof9lhorttJyg2x49/YPIpSO9U3
ZTMGnj4Wxfd1sRduRNUsCqxw7LhSVtgu86oCc3yW1OIqKq4k1wA2YUqlbT0FXvDq
3J9vQQaizQ6IMDt3LA13Thq0JyPYKZCxvkX1q+CLRz0HUyYO+uH/NlNyCQhICH6K
WEVd19EC+3J+/IyF5NTfDLSc8g8tzuz+bdWczr9ies1J+K1LBd9bnWujtabRgFsg
k3Kp9ZTuSmgqo5H8g1vgwOeogfeKmeOfxpJX9Mae4up4uDb0GsMrgvsXHaT6MvMY
9qncQgAT9TkFg2mq6F90itr5NaSHE01sxYsp2jzfIKZK9N1MCQpip2Z6tmzbz+jI
pLZKw54ibysQkDY9xgegL5nA3/rgphxwMsGXe3zyI0KgVUwo4yN200iNC5aSCKzN
xEBfqUB82vRgaKXX391aDOXf2DujWi1CBOjmYo4qarTG4N6h2C0/81jpQci9hcB0
+gg/fmYFUIraBl4RXstGuEHH99eNCXlQZIpUnIg86/j1m56TwweEDvurazECcxM3
ut6ed6mi9GFHs1qyfbw9nTdX37X8WCnrYOIp73MqsNZbt83yLdwrJ5CPprypk3WC
nV72pzjibbobNhlMxoELVVIoDUtie0L35Fcmo6ancinqNoTbK6PtVkJdyxmajP+8
sQTywTTPv3mjXgqNuBmcptRVfMZTffixDkzl6jblSpDeIa0HkuN1SgnXtoCBN86z
mHVaRZ8Qp8A+Rc2gOeRY8r0Uvyb+1msIJnsXvTuynoTMRHfrLinsWP44pm8gevPo
QRUVo/Ye9W7tOz8tBuT2kkVJOxrPPGJNJCGUs/jL85k2Amzb3wF/xntKfLQb2CIU
GgZtiMwnYfPSk6LrQoZo7EkjimQC8gXzJtBJj5guYfEVBYf/z9EsVr/9h4Xuy0gq
R71P5A7ZiiEiZCC0eJs9Ws36i2rL5MXWbmw32kctzTsjgCxcUdCpk/AIHIGr/OLu
WmsXFerObsFQP/DyT6OCLDEewUKtZ0Z1TKeOg72xlIRzJgnEzqHkvOmbCzKhKyUI
ykjNSkRgh9HpDZb0Zu8SHQd/ZC7j60DlQY8/CI2TiZQrj3WP0k1HOPUj5skdz62w
UeS1H4JIXDKEoVip2/2lOQzvy475oQC+jBftzG49Pv9ZIDBhcvr7lj0W4eWkbGXf
fUesN6tzkpVhffq/XPjVgw7go8BDv1iYS/aNhGpq5Vz24Rarkz8b5XX3O9Sye8g9
WkxCfNWktv12gql9sXbdlXOKaqlEz2S972o/rSQ9MYm7Jn4Gb4oL+yYOrhvECqWo
+DYo51q7qo8BuVWZ8a2iOPoXI0A0oe6FT2ZFn68QnbFd+K/IvyFmhMvza/bTO1Q8
2TrU+JuiMiS6tZ50jFxGHfZrUp0z9+JjhMDDHzjkuqOxLVU8imyy6n18uUYVk89c
B3ab+NN40SYuBbBH8OTr7UO8+9/PQcxwIuWeV9bfQ/D+ZuNopRA8hkusp8rHaGV4
/5WgZfe6Fl7KoCSxr09IH0CuDGKiCG78sji0uXZPSZa3VfjVK2FOZ+yGU6BGG4EB
+IqpD++MmP5R0sTtVDcZEtC7JNd750HSOqca6WajG7ZUWHKEl3MVjUvQsYAKk3rG
7+/4TP6LV4goeY6Z+wzwu8G7gfk4WP2cTZ2q4qVYqzATU8lKFLBzcIwrvaY0vY9u
eqzX4DnxvFLz8pmhKtF4MHrITdBzEc6nJgXYxovZmNMMowfe7BmHjyYdytel/YNI
KrKBTl7cvhINesS+88KjyeCJ6UnYxP3I3tuujEQQZYW6ZI0hRMyuzruMakQa37bx
fUnYTlGQ65zmG47o+w7D9T19DaXLA1T1ImHTmokUEaPr067zvd4pUj6lcklI8hNi
7x771msUvEQOVfsWb2p+cipYAceDEg2lMI6i6Rb3Jr1QAny4osYAD5mCTWk2VSkG
UBptKXoejZOk3lp56JYlNx2RIE+hUOg+lxXYi7wBZfYxC4t8oup3FH40qS/erEPz
bO7keo3hA7NTl+vdGTPtWRoL8k35GWQpWBb846QGJEgE8mE0IzOz0vSvSUu5hRUZ
GC8squiJ70ysNmOa+zKJ1M8BHxyCZyuqHJ3d/zIWdtPZ1JlJ2vNaVrzLhF9Zt8Gi
4wwZdGYJhwWoTIUi3QfeH7VGWHg2jszhyjX6nI7rMvNQGkkug/3HqBg8KqzrHT4K
ld5gda3Ab9tXUotxDWMhBK/weKpySYRXdWOByrKXRWR1NlbRBPgBED9eAYNn0avw
1Alk0EIwJtu+nroeCjGwkpgBJLVEyd8TCTjaQtEFmPgGwJOInJABLDj+SqYo5BjO
ES2PJ9P9EPgheCtVoo/wCGWJOgrX8VwWx6EveAWy8tpjSYAhOYhrDOTZ4Jximl0T
n4YAAA9KA2kLNQqvuFKOSJCWPjrulgL+v+5l62dJjAV1KaE+cck79jahxVMh6LJb
YOcgCB7Phpkz+1jvUMmDbMyVR6fH9jmM1Lvl/TfVATaDWF7p5Z/Q53LqDU7M/NwG
ZFCW2bVbtVHCZMFlNqcE+Soe/0s8DQELu/elivMLNINfvwD2zrMA8GChRIboasqb
R8uEQx4XeCzG0tPeRiP3cbbWkn3uKwrFK0l14fC9zwvlJ0v83JNKVDR/CWhYX8xk
Tm6v3sg2oFMJy06r6J9SxtEI2ExTVgKHh0K7hrAdavV/FbvjWGBKD0W6mLg/KVqd
KIQWFBcoEYSg+sKljM51pk7u/3uAeKPr3T+Jy25mFfqA+JVtindPVAorMt28ljqr
bQ74jQZvV46dtBwTbAMR78i6lld41/7sXdSSjKydMfZ6dk8Enxe5cMEaf6JYdZra
T9oJG2M3AvtNk7txC9WOammZA8yoT6ZTgJfIiZB85v9TUTINXtzWpnPskh4fTZvZ
z6pyp4Py68GTQBf66/rxNnEE8OKSN11BYQTHaqtNYVoarkJkJhim4IPlWEvYHIlJ
+RU3vU44/fPCFXaq7sZXeJOQLIbgL6inD+3pdI9M8wqsOV5+++PsoDJ/nDTBroXM
Vue4wQ1ZxSj2sjH5oRGsagq1uy+S+FcCH259EIxMiyOFH33HZmrRjctAOFuuxU2D
FRlhlP3leom6+MK0xIgUcvWaDc/Dx5D5EUm4JHXWfQ1kmd1Hxdqhz0zzPgRVwTbH
YcMB0RtfziwdZ9Z9i/v3Op99R1PeHicY7/EZWBlwczSeNd+X36eNnIQEwjGKNUz8
PqV0DKW9mAhhsvGnvM/AXfZ0DlFGlYTH20EL6nsK3NQzS06JWN353yUAfII4q/QE
X+cR+JY7/DhAinJ+8tr5dVRE41ktWlSEC/BdXd3uAdfeRERfP0yW9usvm78Puptl
tu4arNAzC3fW/NzPXFC4m9FT0sCPNYTUrV9NfUFpQh+QzjzZa//UQBriHgyZNR7I
TZvmsvkW7pbGeF3uWyzy2TJtq4odaZILQp+X2GE6Us4mnEFrS4X/NWySI9jINbDd
PtX8P1xGwtUDnI6UgbelPNOXQlvCRdjMKtagm5hFkt3ezvMQg/kEEzaxT3kw8PW9
ujumpv5Q9q5g+CFp5vOvw2Osnl3t2zX9R9aghJF8eZTvZyc7J1Jd+neuYZGfbq+M
bzN66ZXfVXNv4E5CgBjQ19Rdf62f7ytjC5TtMYrGPvy7tKJW275fvTrTyjcTtfzF
jVayo6v/8VOVOd4/REhqCU0q1QMwKqkveiF7iTDLFdD9sRLbsaW6abExCIo7LugF
MdklacNJ1BuTD8AcEAANeV8I95hxWGRKU/msrSE4KFGU7qMFutXF29Qcw8RbrqDJ
IsheZMVbbI5C9E8uvl0ndM/eSj0coMBqbOJOe1JLAYkmZ18qMLOqOin7FCitWoHV
TsNKZ+K+9nOgWttnIE5xtDNLN5+Y+lb4n6UmqBTK+i6mqkXau4+OD7ArsuEPrBBd
89JyTEqL6DQ2NmkKE3MrFHC3chFBBYxfypMg8D3YTK/BDF2EPpbr0ZHvt2bhY3qi
VEfqx2+unc4Vc96eslBZRZMh+5ZeVkAGY2Dn1hQYc7PXrP2rVAQyXjZimvAw2HVH
t1xmdhLu9fuAADez5F78Qp7cIbliDCsuX5SK1s8MKNfVFL99KKxHfLQkBkE8Y7VB
LCJFW6pc05V9tYTrnkuumjqxkpllP2idUe9Iwlx4i2AljDEKnbTZTdM00FpoEHEU
ch7nCk20OJWwGMuY2IF7l0Ugqt6YQ1lLaDH4f3mpLTwJL7jzTht5X6Tq0Ib+rS1Z
t3yRfaqUA7ffGGuToEfSoMLNiDLEmH360pPx/mL/sFvOCKjOHtyd63Rjim05S+Xe
OWRtLOapYPK4vZsi9KGIKYVyOKXxEmLjwViyqrgY2gLQHgKcktpsjXKDxfVNnSdw
3NU4FhkCbdcbYtdiBH3ZOb3X1amDrkbc1J2gOLnu4vZtLCN2pATom4dFa398TvRr
BLYbRTuv0wBzYODYe9wSa/jDdonIVMO/pQorwSQIarmaJPnxOlBOSv6UYtNezd3t
j3r3p1nyXNwiCQ7g1Tuf8v7gndxSv8Xehmdcg29piXutjcCygXZbmsDdl7FvW0gb
d85vrb84ZhlmatgELIxQBZxFYfsXIiWaJSVxFPvr42PkA9rFHZmnBrn8eWPpOXQ6
FsEhidvkg7A933DszIWnutmg44PWADFCQOL0ak2a6kcbp/c/LbptSrGFXOqwrJTn
9RyjCH/4gbtJ5l6cgHNqE85g+FtRE5usxIa3frlmo01qf42WLcckdRPIfgVSDS8Y
CbU/ZWy4xoGGQG4p7k6MZaW0EizVy9HJmP5pQNCIStvDx806ALfFu7y7wMOoY5qp
skpnFG/JtWg26zi1s7Gw+coWjsNOpg4UxQg/JQux+bYdHcdb2YPhXmZnoBUhUFdD
K1DoTqbYKHw5gZsS5lnXzxv7KsoR7B9MIGjPts/SKasSRuxNyJBzTa0nc3feEenm
y15CqFSEKT62BYT/k+0iHj1S+POaScnMyrZ1p+gL5J9XfleCpWm43vKgRE9xCtNo
s+YVwNSkXYZIXaTYqCYZs6ZAcsXjRPkglT60KRJ7IwW+fe2unHIMA7nb6c2k3t7V
yORnOm13g1Lltqz/4yEbBGX/zcSdl6VN6SivvSpdgZQsbXsxM8Z3i6a9G1qttnjM
BOmAJS7pyZgWmcFYQzkWG4pXwk8fZHbT+JAq4uto6oZhjATwMxJf1hnAhNPm/F27
zVn3iBS5n8BpZQNru6Lxos8VPlR67zc6BtZWj5fWTnCwKuKPtZvzt/QBwxs5NkdI
q6+tihyvXn2htKnWoFk4SJx0Pp3PEr1LXREJIW+hp+plUsvZcr5IPN4mQOhKsKr4
GhWd3xqeq6MnOx/sjKursDecfQII2nODxhoLxPQEx5NyjEtVT+8r43hlm6laEd8X
6uDqn48K5LZqcnINyzjvsemIeCJcrdUE1Kczf9M7djNTRf4SEeVfYR53P3OWUd+7
XfdR7KQ2ntRsC1CK7wTiWdAl912XhzDI+jNM3kQdbJIuq/cQuFptaeHJYU0mOk68
jSusRGZLGs9n3XAjQ8ytY+SftKa0qO8tf89bxenICBXA+RkRsOu4lVc+HB3nm8nW
NBe4SMk1DWhPynoD+8m5J6RCEORaXhL6PclIxR3WMzyDVyc3ol+qylwx/FT8mkRW
EsgjIvpY+zovM4G9WYy4I3CPx+MpGNRJeQBxHT0AJa3pYB5+Gom/Jrc+ffJlXjM/
HLqbl87Sms1ghiWXLcvqTLOSxv53JjLYeNpCb+dsbI3wHe4poD/VZgbyKPVoFHvE
YEB2apk/WTT8u0wr0QodDHGredevizY+HqC0O7UfL52S0lJ6ao1PLm21kP1WZAwN
Qp2kz1YMnSS/FO1D2EIOpQZk7HcOLG+eKfLqOHgx1tiM1+WiRgzwkPGhB4j9LWY1
JNBWCPfwQTvXqMa91vnN40B0quSi2exLNhtPM9RbE9ttYQzYH5Espi+ZfmbRjvhS
fFu0Rz5lkZDqbZa030kw0J4fkmGNNmx/N2m5UO7g/xQXSA/Tx9qF1QpfZPjWMb8i
EplbM9doTAtJF7Fh++fQ7VExpnuStBHj0jfeaLBw8/6DtjUtV6r/6It7yqzV2amH
6ds7noku4H3ciMVVyy4io4iTzHQwlN6uT/nUGdekxlfw37XyifCM2adn6LrjGbZk
ax65yBQ8/IDVrLdTkp9753skTcYVtB2Hc8dzsryLwFlEI1ZlvR7TBkJ2u98fTwr7
j9KGehS7TEQjmIgabfsFRQ2qjPZv7IkrUn2dZ2JbvXVRaxu/9A0wiUE5L4jM1iJJ
wgwwqqy1V2DYawepi6k/wWIsYaNQlQBZxdwKe/nr+JJ7gsvj2YE1ilVSxkypAjX7
NMXK8dHOkdlcZ1kWprlxbxqzrtpQbH0wFqhUuYnN9h6kgHn9VbsBKFct2hSnnRYN
okync1+fCv7L4LGVR7KQhieRZbtBfudyN8wgyNgNWjAA9teBu4P7yqgmP9t1Li4M
WP4h5YNtpUfKIpCj7EmzHcyPMP7NRrxtmLUqZYeWQazXiqqO6kOwtw21VnG17jhp
BPCe787edSWnDZhZKNIzA5LDIv0tlUQJ7weT7AMgipqKlCZq/wMPpPawOX8bwQBn
pGrkyFWxu+kLE/W/y3DuFr2Pd9o4uLdgKxRmakxLgep1SYdubqq9fbCWIIVHVKFi
piVBCTbrT+/8Xg/PclNZjm27ElFYmJURmsG0jCZeHOFAiFTNCBvZO+s7Tlgg8oTz
aiqBGKkPlLv/MwvoCOL8JRMr6JgtMsrHXyszY45TrfSsgLIFT9A/gb6uW/+u521v
8vxQW1hF75VA0Ll6Ig+q28M4uYcCs8PsgJuenJLyiVebIDKkstRyKBXTME5LDRS6
b55KNNKNtPMWpWq3gsLZCAiPH07XpfMDhoc4pBQX292Kgps94Ivf+NOIB5Sz876T
GJXEWzGAWK2BGdgND0BQSjV0UERkkCTW5sqwuDaFZuCD66MfQXrIW+DYDYoQX9R2
AzJuiyzUnYtHnyY58s7UlP/1SLSODkhCvQ2tyu7iva+KVzqR3LljuWCUswxWrTrm
TXwPylvGKJ/mRA76UvVEKfW2/3Gj8tLp+2aRJmQwPnOmb2mz3+cEPKe9J3EFV20B
mRumXEcjUgd+lvhMMj8Mp3d/GRqs1S/pqQPKZpdK/Zb2UlVLppea0dGaCctW0es2
X3ZFeFeQLao0YH/sr8x50lzw+NQJ2RFlMfWRXbFAVvqEg3OIvg45kucv1jOlCN12
lmbauyKrzsjBuWSI8xHVigPU4RCxu8dti5tQxnZCpfI1iN9+j1qi0pB2gR6LMJPy
mOisi0yrQFhIZPhmc97LX/4wPQj3ZpieMwGjlE/m8WaSMBB7FS042g1nQYVo3/dN
Ou5OIhCCendkWe0V7ds/QGKOu+z4mEMeB+iGEb1QUTrVbiXa9GAi28ZZb9nhJTnX
iZwZhfuGK2RnwjqquI2xbUUBYS5tV2MwIBOcqxb25E25sQ8nq5DvlPAhEmrk3KTw
9ltwziU5FVC/dHxn9Vwnt79SJgiaIobJwjv7gMBjH0h79AtUD98MwB14dCCSj67I
jz1UVW1qBs2CTFtoNFq6/G6+2ih2RoiYOoEGIred5WjX1E8gcl4iRXKRbtBrwqSH
daLOMfbKqNw1FLfcXqfQd0nVK0lveWtx67ABizBwXdN1bZXR4zWXROaexAhFfgaH
QwGEs2mM6l6PSm72GnBjTr9rvnqBBKLRhQjzCaNwLjc630eW7SM8JGU9dTfMhew5
OjLVGARAH7k/v0WZK6yr5srT3rZ4J8Zym37Fh10l2WOEAB17FwKgum+0OIDzo5ex
ETNhIQjRjOv79iJd+EPFHAnHDqMbzB9UVR96XSwtxrHrLPD0WlAXYGjh104w2hnz
v4ai6/eIwCmC8t19DaGF67kHyMP4delLnjK9LZMNmV8QnA2KQ5ghMQ6ugtMR3/cT
Rm3C4BqZSDlRdHxY0xxm2lcfGD+K6MYN3aP1KmNOYU43CjnkNiRJbr/i5swXqoRN
8wQZ7DLUPQCJJOdKHhusc+z852TQyX8gOz3q58AO6LqQqg8RHa30CnvTXHSKUaaN
xWY5bCjZ/pRLxAmFN+LGM0L7rzazwd+YVSckil7jJHz+qWBQKRwP5IKcGtAmZH2b
x7E1eRsXJuh4riVZJpIIbpkxNc7tvCn+3QPZwirG5dXILi/yDVctGEX2hnK64hqZ
qyPCrm8W03qRLqbMeqHfXfTTHMGBy7INNmQQCY2LmejI24mjTWTiHZFpgEeiq8EY
K4pGAlGGWGpTv6s8e6+cZveQknCNGuE+TysMISJK8qI/DAK0KOspy2cGyqXdDXe2
H3Zjw5wy95ROVd9KyeK539/mLJLMH9VDuUFt9FM125BqntnMDyr/DU3Yw6Sp9lHT
HOVv76Zv/RkKcwDBKUwxk6hqSIsnfWwSOl5DspwuTaAkTSg8GZyhd123EAwomxit
meLGH2E2MmhwD13C7y/nkAphbVmmeSXjcN6aU1NBdY7N0fYtl823McBMt7cFSXgw
9XE5GZ0jAmjyL2bVb5LP587GSoYN2uUzt2kCM5sKvdGfHJAs/d1VIThyGdqgTEfQ
1KkKX30u5HE1zWVataeLWTqIICJ7FplP/WMDgFKoXlD50YAFVIRz0zerQW6S9PZP
ZlXOXIzXg1KBLfUGQbRPJD1xBaqWOMf9J9f1zP4IvRv0oShsbLTsyTxrJ9HitJA2
cnDgdUK0Qm08ycOXA6lIfeZHzxxT/uMeftRmN7O+ltiNUoTSlMb+ZYQpIfff5uXq
E766UGUggOLYZMRnXiVcloeGi+6TkbmQm5IvpAV6vm6qTQgg7R7chIZOq1a0uWN6
aeiqRFusxMNwrMEJVZdS2FJ9/JDbHYio1z+kskU5XdfpEz9vuzpo3YUkbHqTcX7x
Hi8Xgghz1ZCJeKSkUsImBgE51uUABwHHwdmIjk49MCBhbxMKBdO5ekE3B3Pv6Yzr
IAfXtdb9kLGrZUx6Q/tH7YdoN4R1rLwS7Y9tSYPJGjWPHpeEOcVwPl4E3eWNFcmu
/evgko8uCXRiiGJWYt5M9jzkTDAQIzywKe44FKSx8UBx8iRNgLZO7BuE/mv3UfGh
LkmmlRofc6MX8AKs61cl+5T7PBuqREhKX/6RwkQbkAdKXPIBguIKQf4W7eL6+JDz
xyfXh9TKdt9BMetjvJ2z8U9J15q+uAaO6Z+3Wj4TIgBy/zCc3vOXuX8qAQ7hAMph
oJ0ryFUhU2dI4Am/TdIPGIy6F5cRJTYJ7DOLXB4Pt/HOJlJcg/oLXeeBouvO8NLR
4F5e/XdNlfQfdj8tSgtyJEG/2ZARlAyodMKp4MmYe35M49OWggWVqZrg5fug2j8f
RHmU/K79OEEexaA7EwgKl+CJrNGbjMs0WK/ktuaTEoaiJpa2u6RKd39uyKULd1DW
6XH3R2rUdZYlzmm9gdH09gTywZnjrlNI7xgMY6kefUZZF2jJVXWGJZoUsg+YBw6k
24de+OZ72v+FMYLWGTGZoPcaaSC1gPqd586DvDA0q6rOp6Jl7Adddu2j+lYgGqLj
dEaR1CEhunfofwlaSNB6/p7Ek4m4m76QUzbtS3JC9hKw3echxABkuZnFWl2YDr4X
jJFMWW6vXaoZ8ZgVOAqSDh9Yt98cm4FQCbc0Uz4CxgFbcVlUL/MVWSHy3sd9KCdF
lOg7meutZ18qaPt1vmiICFTC8wKB1NREf9ge2NVIQ4YrJAIF7NiGMAL4BJAueNM3
ch8xs2xffn5sFvs0MNd/RWL8XXYQwThLdJKkxz5DegW73MBKTiAM/XpbPbMFqGYk
xXxZncE3U72t0E3x6ovDD5JNEPMMxYopII9k6hij9wjcsrvUi0McaXrordGBgU+J
Be8Zo2wXu+iRny1QtTl062r9DDD4P+XO5pJibshqCdwPnyfoRwYJIBOKZvewivxV
ouuSXtJ4MFydiHKs2Ab12i+DEEhtK9VGOmuYLXwIUcIkkab+KMP32chkXfZ9b36Y
IsUI9j7RZR7lV+2xQXVK1oidrA1WGhi/P9V68fqWjmvISremph44r1MC7t3P2XA5
yLfcre55yArZNyoPoI/HL9ju4Ru//JWbYVzNPhEU0hRubz8oyAqKyfKg9UqP4u3C
/FYfVUHGxgGJPpHZKos6//532VuaMCx5sUET6m9aqoK44ddL3WLoPs3fIWc4Y0TQ
x52x9NlIhXddKVrI+O7+/hVGZW8Ekj+jexlyxEYUU2LrlpPk2se8BfiQsHTCIscz
S2BzmOdc2liteZvOgkQjgt1EkN0rs+QyBaDX5PTeMOK1LtzjB4fa7Fehiy9D61xl
/IfLlKc6YSokr7HrBYe6ss2C+7AJmiaPnk4IQO784XGVXZl+WqIDxm3zV2JZQpOs
rPOb1lJSnJC8vubMeqLySVYzo9rFnPAOUOinwEhojEcws7aQZ0dcRV+2CaMxBhXs
tI8NHEsH7+cqPc6dl4vkz562HoUivN8pM4KAYzJhZDE36FWujp0BukkjekXtdUNH
u8E5tGqLf0pd6HT1kyahztKzmAq9cr8lkzeRep6MSC7DrRTxGhZOczruiCrLMlo0
shmhKrnGxgP5l6aueeZI1s9Fjj/9wdnqA1Ex0tQo8d81BqnM+KfGcvscesXQdX1l
UE9YDfeJs5ZzkG2UhNewm/GLAQ4pCRyY4Ryz8/UwIPL4vRvEEhXras/aUjeUhT3k
FihkyFfdWlcAXCXMvRngbFWNzdxMq8TgYwR0ZI/mVIF5VLshZ1f07Vl9QRtVGSUd
bXEaKeA5L06RWBulK/eiIuPEhupDubd09W/Ltg2//jb1L+sY8zK8BYvGtQ21eFG+
XP0vpg7JX3wR6o12KirnneeprqhJ76XNqGKOCBo+e5fJKah11pFoD4Nkwz1DsjYu
v5wCMa2WWvSgkYR8sUcMraPQFkh32ayGLv1s4h9jRFCDlsc66DXRFHaS4AKgoxF2
sZ1hGEYkjgtmETRZQvB675t8dpX2T02ZZ7FN4jW6QNnB8NLKYw8oBafXB4G+cFpk
wlxQi0F+JlSlwXvtN06T+D3AWWXPRhpAtS72X03zMbreOhrKlMwu9e40a4UOxEqE
kpgpwkpxPucivEWMp0Ux6wJbH7RISlLVhR7a3DeqO22Fzq81pcgfpa5cLD44Kjmo
jxJaTeWP629hfZ/AXk8RqNUcQfM7q1zsJidBwvPWxFKZm0O+Nq8hMmrkL1ipbyrd
l/s+k1EbY6h2sOeKkyqEdfKr4QVUoAs9/26G38ahyRB/T/9KC+i7zHtD7NPG9pmu
b/Em2JYV/DTjd9AMqC1RnvfgKuBwj0dgjO06aqo4ViXjxhmrVVQ6hY1GgMihc+n5
iDcS/q2kw5bmIaPsm30QSROcr0hnKD0MQlY5Z1k/qio2Nn/q+MMeB3ft4YQJ5tQU
QUS+d3/NSaDqtF1NYdxW4i9yTfIJlJSg+NDsfE6TBNiWOs0f+3NYUSE/DWntnwUX
v38JOwkOrclMASc62s163q4LmICRHj1CCTWsvsCaJDaDIB6d76Btn/Xz35bZjfJb
uhEXVcqdQfXK6gz06YzMIt7CjlwRjexfNiVkrHLQw9TN0U8GWrIWj2Pc7YjyH7k+
iCHQ4bkGIA1PaBpDs8fGnOekQJXNIWSztwQlHAkyhriscQ/HBvuRueKFXm3V/Tk0
hy2GoiuzvJYbwxaJz3FDfhfsKorRI66/vPQWPszccrA0L57nmiFUyoaVyKOwYq3A
QKJ8zczAEEAKr/98EySv/D1L4r72VSDnrBgnCNtdGNrcSVvRYc1fHRYCZ23rnf7/
/tvUoA876KjbGznhndMtEyBUvisGgf/zyuUkfbYi5TM1Z+VyaWm390dWkMLf4c3n
FCa9fjiHLQz98j7QBA5wpXORD77Sslsp3E717R9F5KcvcXSugiLldGKryTVJg1L0
/RbOP2xBo/OygMObBqHWsKq8Y0+DBwhDTDfhb9wNTidppfhEv6xZP8gPBFxBl95F
wjkeLfRGr2QhJtiH0y+a680Aa2MsuZLirMl+NyvjAQtjNau5u5TShDX7Mqw0v9+A
8uZTXhlbYc+shTNld6M+Iaa113oxuTw9qB0+oCz873QlGCnLYCgy2Qkv1fVx4OLw
Gt6xFrHWu/QkZFBxMH1lsUf5WhJiqtnWy9CufIU2z5fwCz2sCYm5uar5q1XjdAPp
U1zq0nbAAGipvi5csmd4apq+BYpQ/roZD+a1YjMoiXBwKMNlSiV/tM7GDgWMRoyn
iAgohc+u0tUSAR/TVFKBzlxd/MfAm/1hF6zCkuHoMze410MLEoVK1dVIcC5Xq6pw
Xr3Epprpij48Msp6VxKAyB43MDNnXZL/KoOGWqAPwvWMSt5Kkj3UcKuGrLFyduQp
VkQAPUqW9nl9TDSXSNnJ/JtE6NGoDFEbC6AE2pdlG+KiVdz+DnzbZsFRNJpIX/5R
SbozxVv0QQ5XvLYD6SPbZn3Vy0m6sQJl4+wDwINWzV6ZbCRASDC0oMNKpyhCbE/5
UVSbTrvdQ+GUAWi6jV6QOk7zg1XlsV8nQ+MccfPxjUtR51p10pCN7rORxu2AqQxb
Ujv8qfQMl+kpO1TAQvncNsjajQZeYRR3p0x5y0ZR82xvxyTEP0K8Z7KdQf1rrjqU
WGIrd+1XahGWQ3M0Ck+AnmCy5p1q3FfPttGg7KXmQOAwaC3XIXtPR7/691W5uvvh
6Gb6lexckQN5yOrqxIzpFViZsiruJhhz/60sxtVHpaYC+8XPUs9+EWJ4q1T1ox3S
gibqa1AkaqzownCctdqSrmwKQGn9cuHW4nb9M31df7EQEni75YbJSZYQXjOxXySM
s7aTkdtXi1I/jvd0FEWkoQ4Tuot0V2FAFztMDM8r+hJE9HbclOtJtXyOiAMuclid
ISXzRzZAjeL8ugOKwRpae1Vl5TsforgpCiK/48mgFE8V60qemXm3FIu4Kyknl8zx
S+heQQByW9D/9DJ79d6egPr9MFaQJ6AP12DQK+8JZyzIPXFUsmX14Jej7mvbjxT7
BXvBXxyW0Zttz10g+Sq92R7s+tk6e2rag6jC3o3nlLYF1tyLlHbVlTjHTLk1xu3I
/yoc48W6VE7qjuMPdvYPlpdBIj66TAN+Dx7tYr/rTFtGXEHJzcGV8borfn5zGCw6
+4GOIjuGtkPjQ9dAJxuI13fmmiL5aQ8bipXjsE38t4+v8y7sT+lK34zHPW9w0l3W
/Xux6KaAP3r1FTpr7yV6s1WKphrUvDm2R+wfBznuhhf4fQTVCh2+tzbWYwc2pm8j
RYeVUGGnKDAz7FLYiqTlucAXVK0NecR2g43ef+eswBH8N5/0eSe2cGRD6KscGDol
ffnG8w8GeKk83Nz33Mbfcmwv4vUQEboVE2LVWtvkuqEENm1UCW7e/Ppa0MEkvUcR
yEmzqnUoTXtEklXrWYKPAcSvcUZzAEOz6CtctQEzz8X1ZtzOJ8KcuCRs1Xf4tWEt
3pg5m6mkyGdZP5IXuP3vZlmCNLEsQApIaQ1jDZM5UHNjWh6HsM24rNxaLzvFIflG
+q0xUMscwJXsGj6dOv2O3LBPqv+zRRlmzRMMRQHUZ2kaa9Eeyqo5LXCIRywzep7R
o4vbJNfY+xlI6LnMr2kd+i8/90lxtX0qAAzSb4QG53i8Q/GvrzNnY67QJeuzTaGp
oDsEbzUspOr58+utvNY7/aN/8ufpLqnjb2ChWDHWRslg+dPaomYfZkcdi3xt7Rm4
/jiTmj3jebUWBNQM93U6M9arZjFgIZ/LQmrYNjlrvf0cOyUGwkZxh2hsELg9pyir
uVRMLKSyYZJVBzrmk8ECx0wkPJ8j6vFI8da19moGmpTu30XAL09Z9vFd25mvXZNf
qrlWNHBAPV0tCkuAB75ZjGWzwsCExOm+iMFDevSIfOXgp2aCyUp11+OPKLYNGPLs
13yqtLMS5Q5InB9sB8tKfAgeKZMbhiZRBls0XnWXGYiM3OKiiwe79OooRgPYdKhA
KeXAm9H3cWe95ViiHqKTbIchhshpS8Z/o2zPCl4oGNwrFz13eQWKY9KhN9XGqk9E
FzCIyl3VWOtPpesJPtCg+9B/7PdbqDnnKGFA+xulC9JEssKww0JAVL7E3Bnh+GHv
8SttrElxDnklCg8ihFG8wYmkcoGbAOuEs3cX3/RXrWEqjHbE6YIDKkV3rhF3PItA
zOThPe+10BnOoNCU1HVqhqwu+pwNyiK6Ugaoe7aEFxeAbOpxLmJW6D4YnASzXJel
qEiHZE6Wsh67sQVLmLkcaWL05gLPsKdU8B7Xqh5FP+0xYdX8jZx7sa0GAV+s5QA1
qa8QTzMYV0JNL2Iibut6J/x571c9IiL2AjMVMXjGJEWpj6FiHyevB0vvBO5TAB9w
+/WAbubtOGmL0WVUQbThdtzdSaYHlLnsoCeKtbtQFr03iwFW6r8u0u8uO/YToXPQ
5+z8x/wcRcNgp+2FOOGEtoU5SFXAprg8oR3iMOCEhu3YoUkSznzXrxa7gUV++gbu
NmXzutAY231Y6gj1qgukfRe2vB7/D082wJ0hvAuPPn1DpMjYbOZULlVlaoDvoETq
ydznkfhPMONy7h43juJEfkdCPkpEKncMhWK3lUjVeH40hUE5bzHZc9icjJAB3Xfo
IzGn2c2YeYeWV/QcJNKYlGA7J82Vru4VmuNxKxcU8COll585h+zN03+MQ6PBSJOs
087XzWZNKEIt5YEM8v3+oWF91vyhRIKExDxACeGXvNAx2jtYiQ9uxNerPbeZ6o19
2SqBRvHtLyYlWr9sWEmAPIMgb7EIWyyHC3xTGm5B7Jhu9mC52Eqrp65IGImKqnD0
nEEdijYF5PsqldrcpqsvEKN2tNp+Brnq165hcuQj8lFl8wrduAWoCGGtmURFSn64
15hfsmAE6CC5z/yPALtNCGlDZBm5uzxvhF96xsK1CM/3Cmcu2IMiDeTMHEHYwk2H
7NQtzHRIpxzZ5BWsCR4p9/IsTWBuZFeikel/W38/ldBACaiIi6OHTo6TjW5Y4zUO
IOsbMOp/fvpjKk2nZmqVw7lSKBcoBA4LRMEZcFL1gLCnejM0Z1RvVh3AjxydQk9p
GacWk8ORPh64ZHebXGHSxmURRNwsLsuM2U7Ys0KyXZkQn0G6NRWhTRyKWQA9wmtC
7DRenM7DoVbqTvKorQtW1t7uEDN3tPiDHA/i4kYTalBlHkQAGmmuaTdYMxtQ7E/x
vh1mB+Tg6lzjfYww/nYJSQLVVDLJFdVicxTJ7/uWRoYnns/EDKoG8TsYK0bwelWP
6wxC6iXy+Z1UzZWgOoDGETBd7pC1XqPPR/3WxzEvpb9MOHojJNbw2tfbsFlteyqm
d3DXzb3eu2753QaR5EhCoOOu0LVBKi8cLSsJks3SPxFrrP7qcVKKS8SGy069vcQ3
+vclLezosVZQG1YMJd6yxhCHuCRIKGoqo4gTycsODQPARgCSxidoW3gYY6pTPskH
/JbfXkzsuIKB4S8bu0dBzQvXBLZ59za29iTRlYZHWs3/PrpcBGbq0i4VI7v1zQp7
6Rr89KBgYu3SJO8A5oL5ZqZ+V1PM24vbJekbSUBFzoMkr6y28cyTARAWB+7D8DOS
XsnRvd02VjkJ43dG6h3aJs3z/LCbqaNSt3X18dHvkTUW2AiA1DJEI1wwKrlx8OfB
xdtUSiF7L3hAT4YGzATpAR01AP5cgTT2PpCqd2fXCFMa0IkgLpP9nkaAG3tWu1pY
+RiaVYu/K2t79vVH8j5DmarD0DSsZbkkVBm8hVfLLEK3kXZgEtBdsOEJhASx60H5
v1hIgyoI2bQU0IAGbfbrtXx0jLTV85bkjrf9WsmAaXlVqQsUuYGtH9+qus1joksx
kUBSRVfsVjpbgn9fNggdVVGGwXAiMjYreCp/7POGiTAfixJ9B7jpDm8T/ZGwkJO9
/77GA3kOOHzqa+SKPMSC31DuKSz0hlRnUWz3OXd/036FSzyGN6Sa7clVHGfnH8Eq
Ov6wQrDTm5fOj36sKsVFj8iI9AngF+VAEenmPAzsizcjpSsmHbCgKfDt85KdD40T
DIMAVT7iN1ArGk7ZL7OrnWwg3+p8ZeQ/s+az1VDEv8JAjYhLDut4MEYZN1cRXi1f
5sZS3Cf/HXRcdMKgCzVOcc1eM8dbAEFs0l9pKFxRHL3AS4OpNpODPP2+XtY76rVS
XP0hyb/OdDgKrlgiBaZPWugelspgKMn41FBOXYMVTVfOhV/wbUjtZCiIbPFzAZ9Y
C9GWloXxPqUSxrdMjTf6ewyLqYtyHI++iLCe0z4mnSCXzet+hMeDOrs7tM9dgHyR
wed/3BTIdJuy5/IPyKuM7A6eBw4Qvn61SoD7RJonL0wEJNHwF0eqJaF5KYcJBU+J
nHT1zrxBe88y7br2OFhqq/IAhtMos6GbeoeDwXDvrPa9kL8ogu96YQe2A4fTHc9A
pcMEIxVwVdgxqR+90hlDQBfU9NwrqmUcTDeqmFnPLoxMLYtdD0YPmOYU8pzzFWL+
t5cLunjs0OVNwzm3s9FITD/Bl5b7XcrkcfgBH0rf42j6/XNzWtbslwNEjG/tqvOW
/YNHzAn4T0M9joRwvrIlWTX03PqzaumsuVqLi0Eu1ak/EEbkdsqbtIfxIpgaSJ+P
QTbEf6dTSz5xZXaFWS40fMu6wFuFunn85eLBdrccrVwbaZUBdEqou834Q0kSSAsV
Wb1iDlX9EgM8xcd16qGOYHji489dx+sC6/Fd6m4zLdeJtssmhxSAoQO2Rt52EpB0
yW5VuZnd/wHju0sW4yUJNORExsgcQNXcB/c1twbohrB7JxUu3CcW3/9eeZZ5GBHv
A5twlcCgujpp0MZ3LKmSnPoD3JJ6CxC+ubKN7h84qUS1ezqbMctbX3CtPTZe6pgQ
LmyE7+rncWL39hkWf21dLxv8xQqG/3Gs7uIsF8uk2Oq2Gz2NiCuxpsHOsR+qzfr5
4sefR9+7u2PswA5J7iOpBaIJ9Q2M8gLd4Tb6DBtah6X2jY/ymjyW2D2vJHazGs0o
qScDlkJ+gjyQJ4nLVckHMVL9+WOZQLyWe3SD51bjA6zXNov3XAoOKLd+x29UGMId
zLF2gF1AzAbZcENEvdF0tHfNvtU0YrkrzigUaqnu1AJ9Xm+wROnxHfpTVWJeZlAF
5MSzRZXQEeBNRJPtXerY1veDvKy5K6Huu4LRZZjcGPN4g3s2hki426jfhE/ne/JM
itEE+Cn4iMJ+61f+1ongDa01sBvdne4ktHjsmRX1wITJ5NLGzZ0tcCf/SVShfglP
Upf2Rb1lZPO0+xbXVihzJtpqwDbx19gEAyB3kzuOG4hDA1bspfoG0OxqZYVbSOom
9z9ocxBW2RgER6jmWOJHMvytemxKKyb1bVJbM0hEAaJgS7fEVmDgbQg0CfdQikXu
gNZIxiLhkS7CcVjV/qCAKtflb0CdcitDRqZXZy8JKWDcjiYMPWZLjdO//laUMLAf
QEnqSRHhgQHIgYwo7ZlwgI4ywhe4+3uWEa8RICPNeW85TFn3YsLEm0efWG5DSpKj
+mLoj0TfcWcPRgOUDUs1yDkDov/xrfvvv4YKBXlMJ5sKqQfdac9+psfN8bJvRkRl
vrrNNpKzZ+LIegWbNXK+/4gYBAV7Y5x8HFGHUAq1yx4fBUzDvG+EE8qdWQNszlcp
6SfdLRanfXv+w3hhitsVQYn4lC5snZ4CA3m9+oIlWYA2ktiHRyS+JeWsneYjWm+D
W/5KaBKvWTuWFmCVCbrm0SD2O+AqAKA2E+SNKaHD494VaTX5OxOSf5qkyQl68SB4
z5yceBkzxz1NNtqezoRczD9x7DiF+IYMcUwPK55Uq4L168tJbOHFN4nDmDzrf9Qz
d/3LTmFchw2ZzwZbEbGUmJYScnMWZesnodbxUTBPpWyXQk8cCjjn63cgaB8JbtN/
ydzNBCKcihpgGfMPS3WfaZWyiRa/yaN6Zrl1kyPvtNGECF2HxWydxH1I5UipaX4A
CjWjD0rOr+JYxZ4aNo79C0lYlAfLKlWEndcjE5/FnDKmEBCDpY5+SgiGPFQEmzvn
xWcktmMZDNMi7uQFzFkCp0uY7HHOEyn9Bb547WNaPHgdaZEvci/0ktjCFvjg+klK
TlrbOfhjbSNLDDa4Jdszw59H+RxyE5GiaHdM/SXwgw8F8nAaG3SxD24OiUbdzuuj
3KiUXpM1VlqHN9PbWwoObgN1gycgSt5NMtm5C77K3ft+kv2XxHaLKPZ7Zu3W6p6I
N6bAx83AHRjRCVFtPK2uVDTMVq3HqIb+Y+lBNw6oSUvf/2GeD/Br+f1jnIGvgwhj
cbgoguxX9wYrJ3EPQsf5sMM1jd0qSHdkCv1WcvPwahlx1Ex4VCcysBbVRvHm52eI
mOtpeeMrgyhw911+O9+DipZdfNFXRE99bNYSAWJGJ+1yzjWK2+2owle6yFFe0WE3
Au5Y1+Qie7PqTlmNtIune/MqJ+t73eWoiMg7+FdiPNRu6cUq3xR5WTFknAucSnuT
CwET2sxeJDWEzNPPcwDw0eVnMSaiGgyqPTPwh6PlLCi3YU5aQ1/brnzCkfcS3ToP
c3amXiTMH/w8Dao8WJ40j/cF9xh88Wtg6KKSED+xz7ikSmPFI8f64O8ABvp9kU6b
JW4c7/wWqiF0TrlBXy8okEuawQ4skk72ZvFuhWbHFLsGe85NbWD+X0yQGrplCgLT
uG6IBo7IAgfMiucIf8JKwcG1y9X0pRCtsfNytCnw92wz71j6In5g90N8lC44ZzwP
GjRhKayvO7MoTyxaN0g/+/owYlaJLJJslnyBgfF/s7XM5V8wTKRt9EOZiL/JNA05
aDZ3EEV/kiimZCf+ADPV2lSQw1Z6/sgHUHWAYtA5wEai7KU2IEcixDNnU7WWl1nw
lVx1AnJHAiGZqnDcT9yMn9G/jDC6RohYEmTi3WZABII3mjsT5BjlVQmE+lYTMah7
2ZmNfaxb8Ay0NmlJzriYPK/f3XQYaP6jV6BPTog7PgAoFsoRJtQ/jEElv6eM+wRx
LiS0WGGx96USE1TOwJfemCUzjkjYFH0crBdl2SbvdtSE52mioxrRDnse/TEXoAwP
PT7EiTw+z3kz/tw4N84v03Je0mp6VHXhcb2dOzK5lfBmDtjJfyRzeXAoEouLE5RI
VKHXgkZLzdfU0oQzbe/ErElWX9YwcIC4kOpkxt4vfxSKseL4boxaxikEJjuONrWc
Dp/QGSM48mMgTDBGSYKUD0xjiE42KNtQaU34eRxzbGbrvDgvidN1GDNCeGSlLlDx
FBGAwt7I9ZSycVBJPORinmx7aY9FdOo8CwsOTD8rhUHCPGlPpmQDjdW+81yjhzun
8tp1XJRMN5qsMsnuiC/HaH5icP+zzULcvPsHnElBZKOJt55EbtyZ2JZ9mdV6dc4R
LBF3KCbfCttKA405cMckziG5Ap4MAikzmIfe94V0Cfzr2FRclNzF1TjvHdEv34TJ
Rf2UfiFCLMWfA6HVrm9l284InTKVGHXfh0Im+AwtXpepai3LeHdREtKqnxBLM/PK
wsdKPHwXZKQuU0kZbWg4Pxp+2FzB41UQZ/UDl4igDqfl7bMfEOIQ6Fec7aifs3LW
as4Y7IqKd1kLaquOr17o1GFcEc4HG5hMEkh2/ECd1vRIoZAGC5SwsJc2TGbHVTmU
GidTHgXVghTPDLKu+WlRuLmin0GVrxRc6C9IUxoUwm0FWO9aZ9ScHaPK/V2tnTVB
FLi449fCvaV+dSi0uRbeTKsgJX6NqHYrMHEe8t1NBCZW4DlUXndq0t9xtxnxfQ0R
Y67SOcuLOQzNHLA4t1q3hLllXqrGZ2nzDeV9rPj4ulEnY1ASQtwPm/ptcWT9qlPj
IzixuwICjL9wkS3IYWTqE7JUjZS4hoQkp1BKeqbrRWoE0YEupF8HnbUrlAOPbOPV
gsLhQt31dhoHs6xJ/wlREWp4dbJ9ZwX7p2/EgOND650LWaeNqvrVTaFmsg/9P5cA
Na9uTRzravqsbxqwaRJD1rYUzY/kp6bEVEaCdvm/1bgkHeX1WXChHv9DFfeexDao
ZfbtNDAfLjkKHkE3hy0nt8e5W8tRH0Yemlljy8rRaIalI3dMIHYE0f/ohPucuepn
sYaUm+lwuIhyAI7/zMj/nap8WsNsyRUAsIYD/QxY8jjVHJpKi5lH8JsFAg8GgFzM
N3cHvJZ9IVPGUcu7K0aEzFdXish4Pnl6DUh7gKwdq7js041iTI4Z7dwvcKbk92og
/X8nznN6/3Dws5DYySjQd5olCTg3UIlsLO74jo1T30A08i2MXiF+BmlW/wx47nka
oGyQoUxTekPvZJoobpQ9VrupGFvtnrOrSGY5HYz1J0Dklf6ZT3FZKDes5Kv5o9Jh
BXSRcyeChH1j+J1QnxHmby5UrmPoMlbI4boWrqjlmO8A5bUFDPiQdfJD5z2GbzIi
0uqnqTJ2zVj2vq5Lm/f0U+LmEPsuCicCprg/hjo9tTCgTUTu/XcR9Y20R1mhx490
bOOW4m6ub5LsGXphNTQ8cPtbvUrd/NOVsZApihi0z8uX9zhfqp9NVaNmCi60elSL
AxwnDzFyHd/HPPJK8oBNtQ/nyd7bvVWtwd/yOItwNp7PYmcKBrYsvwXtV+bizjpC
oQEI4HSaJ2mD9Cti5i7kENJuIJ/xEzd8KQldpGDDQPZCCOHb771BNH1qpWZE106o
Z6obs+wG5Uhiv3LR5q8U/GRais9AXolxB2TkZ6vtmJwUBn9GepKfwWTb8mZqabuI
4QrsZpHhNWFCOq6VLAg+af8eqF7Qdacpeas3oANG7fhU76mWkmbZKhDk0LC5Q9E+
Y++vZmD1whdziPON+FGhoV7/Cp6haQE+OjAPDq0QTfPMZMGUi+ZoblpF4hSwCYOE
lx5R2MglmQj5ZIcMLp18dV950YzOACK0kj+KqXb7k9gHAj5biVywlUspvAS8Bjo4
m+DYfmUT3TQuathwG0qU2VdUI17kP9x9ArKX2SlQU/BVj98uvdJQgE3pSADXhnSX
6Smhg8QDo4C8m1mjudRigbo1a8wk+RbsyZmoIWDBKCKDKMxvfqUT4hCtQvvao25P
HhGwS5zETwNCPgz65sJsxT4Yzoo/NlLv8EitV0CM45LFuu8xcEjdvkGziHvexpXG
dPpWBaSPemlxpMpTDDYNOlUD8RWdukqbipT/f1iOpT1hhMjWM1VVI6dnq8ricU3T
ipjOZt0fRaU1+JcWGO8piNSWlfnx/8J2fXa3R5PFXu4FnwhldAkRgEh+pBlPHrmD
cfbeYtPFE9tRHfKCTlTSv7eZPsbwpc5aANPdoeefmdQcppfKS1OssmOD9j+xb96o
ggtqDzqrhWE+S5AqE10yvhalQEx5qzFM6NKhIXh4OYIDnMWOssmkYyvFDA19OG10
MEUgpfHMq9OYTrIHgx1+VrmdDEl22OgqyNagD3nlnN3Jnszh+5FOFVpexja5Lote
t24SGHrrcbY7Okdzq8zH89xuL9GHsL0d3xNZke9hSk927hQzXfit8rV2Tj2e1WgX
LmAuqEw0xGHYeqMqneLW1O4P7f2zN6dRi70lYlrP46w/8MEdK9Aho6DDSc7ugiV/
2NqnkTpcC/d94/clfinWrFEZSMILO3iDGrA4tYaJnkdlag4hhqjhyZ+pr1adkVIp
QCWFDI3GmvtanNac+1IEJuT6TzbPKm6ceYUduLa19Sh4z+3cO8AlBw9TK/+M73y7
0Ng3Hw6KRzpG+ydlEhtKBTa22hoplS5yJCrQY/1N9hhOtd7X2qq+3kM1CWV5T2gK
n4eG9AITiI18rvJtxSSOklY6ykuk+br9xTgcrBvSWftm3bnRhxTvmuLmES1XP3I6
nXhu+jsY2y82eqYWOoL0rxjcNhYEYAI9BlKHoyXDZjO00nlj//cZ/EHFnQ/BCMlL
RYEvZE2UuV1//kXGObzwUrFp8bbluhA4T4g5Qa/5UJ1M4tUlYXL/YC8iq+4/1/i/
ycvyp1mHsg/SevcD0ZMiNslJZJRbX04t0rgPPgyTu4UAj86twWV5okfgZvZv5D7o
rppsnnU+7/1qNgyncfHK0ha19pW4B4zlVNyWMKVnafewL+rURSzFB+Nk3T72DDWD
3A4k3rmVJHdXxy8BouJyouiHybecA3PwsJsQcqYFLVfGmVz75f6IGhNLf7j15oA5
jEjRQHbmWWokTn4twsyASEwKxAwrbIVyr0afrpUYUYXkXDhosU4QRBkZKxZENEqM
JFcbFO2AvjarRM1DgKL91PTjpcdcfZ350wrs82bw+wTS3nI1d+75MwrCkjfIiZ/m
XRc1dv/jWHL2B/DmL2aXf7zjBITxTqt0B/2Q56PfRi9qEqFoVNk9yZxpocZhgBRg
7jFqEHt8uuHVvApBeAeZVOnr/dHEqQqllSEUWXkntrRQe1k23OWoGAmmbb3yIQ5F
sErTGijm+E/df46aDL0gAFplNIkSLwwFClPLgxmX5K32sWp/H+ZgRUTbAt9D4n76
9xfEoIlA8vMTkXmUo18PlTN2eiHxt42ynbeYFT8xXxDacEk8BkxNWDQG1ia+O4+N
HZe0oSCP6cEIrc+I1hrrUI9bXIRZ7dxgcOhDNwLCpAosjWQ4itXg75s2MovRe2ug
uyWeLS3JRoAf7G9CKQx9vPis8eH+I6q/9NvDKyDJc3YgXi/gPwVrcgL2NY7agAsz
Vhm7n+2yMQmJBxylxNeJTKDx41fhKSy3/bjfL6FjMP3Ral9n4jCr2CN/nMuywVPq
ZgR30UHc3ft9QcaSzkKNaanFzk4EiAXS3wfO7NdFr5s9StSuF3GMY0p8IEh0XTd8
3GEp2FEbIrsK2h7hhC1+ZEp3Wt2YqpyZB3IfSyy9zLxD8dRnBD7TYQgcSmRvZnoa
XrjyR7ES19LjKDRmYLfsdbxsIA6awYykDpD0cqfRPGaaB4he1WDans5ctfszKabl
1EtMimSyzDX4qm6pzCzc/6U55ABzVmefP57lTJbEnzmIBL/xqeE59vBUeo3LoAb6
b9sW4cTjvsfr536VoHctzItEIFpI8Yb/cBX5xXKCNI6XoUU8XPYFtqepWbXdMQhl
v8bBYZnDsSkSIJTVQFg3o22Hx8/wazpk/euBPtgUHT7e1m2cMspPRx15GJ57bZD+
dfwTABapRraKWzW4mAx3MtQfvOeXLYBATGY84NSTSAYRfO8/VLDZ6cyj85xgeqXj
DBFONkXMx7p0qykV1gALcMXQUHOCZ1YMdRSsTHchVf/oisl/qxF6X35n/v/bOopK
lUsjJEC4PK+9H105w956XC5Jt//rc/SMnhvUivVwxYtU0JQYiGz4DBBeH+avIM6L
cG87bI7bZ5sDV52BL6F6J0YgJYAuwre1v9kMiWNDNwx+luI7LNxiZW201H1LeZ4C
dSHutI0uaw9GvgnnneISnMVKIhAib3ADbd+u/R2FwgRdxVRu8BquTy70vGwX6Hz9
jwPVZ50+m0yylVbxFkTfuxfUwO9+zlFm5UnkTpf7Xgtfn/0ehcD2sFoyjVi9HZPp
xCFLjli8GNjMu0CkSNQsqZDyf9qAiz/u2VdN/PROJABmDz3Ey/+6lSSx1kSGUWCI
wy4Q8QufOXGerw55F00ETKcq3JYrTsTMmc0TWfWBM50/O/LRvrmExsAffTL1XR6n
qqN67bKyITovx19mSYBMNMdzorqS7avBabxdWOtRGKpTnFGjLt79MF+SISu439Eq
qlke8y7eZmFf7PIxZw7KOlBmGFx5XtZH3fq/k/L2lezGfBxRLeRCRYfJ5tuQfyJU
OQT1vy0a7nH1dLd3Yw4qCNYVR+cp72bfFofkk5aAiAsv3Zf1hBeJoCOPAOTXxONe
6NlisYNXSEZLhTCdcMqquaSawdhjGLbpSCp+rAir4UNuMLlcKcnveo3BYuvc+qam
6MCSrOzIHOLa/80+UPZOfwY3B3lb4P7m9kBNom0/Xe9Q05sOXm260PfhaUTgx64K
n/WUwSMdyRlzHr9DUcZECLcFf0XDv/KD8UF+/h2dnhaD0fui/I5rhC0hsnZm5AXW
Dbm1vULB5E6U8TxyPxGbPLn0cSNDgXy1lfpf0ncOu2U1hZwR5dajegXoswcwiMKm
mPoJGCABqYIc+UMaseF59orwZ+BDd2B1dF7FGMxAKiK0JWgZ8nsXBXSAlKJlikjL
teaPQItf2SxvjcMpFGxYE1UIJ4woRa/vbjMfb6ekMonAdqddW7MNwnshwVqdxUQ4
/QuDle/9wqibpZMjknxUE/wfw+9Q44jHOOBwde7VbsgUzKj7XuR2sMyPUVlYf3XO
ZOMwYezMTWVo9clC4mui9o5OGQ3zS3NY75HfJkzxyxoqZItD0euSQf82bZavwMEq
ICYwDQSjZLX/9OxFZzzHtdCzcPvPztk44QQKQoyleP/TId6ayXTuUKraNU5dXctr
kZjKH1v1tGFdgmPgE9sFwe4ts9GeC1CW78dz6BOa9tfwuSDgsBRjRT4r4Ap0bJ9w
lQA58jIJKgRa6V0fk6eHuv6ieNX0DZ8Gzvg+oN1ZdEfwNaXkazHg6Zy/1pr5OgU3
LqVb+oyd1DFguuO+PoRe5ARygtzxzoRUY7FEcrT3iADLmKPFW1e0Sw0lnipM2AVd
vGmG+UreC7Shp5NYBHzxHFLP+aLR91XBnEQuRTxCOuEphZoPP8hpmXivpTLjBG4B
NkNcXzgHNSRmvcV+1hkrncboyWHfQV3G8z+p7yfAnXTp90VSuHdJ6yDIMKgBUVrC
jJ/tv0XaPMZWI/sUKuzlgoycQ79ximIm/+N6CPhOMjycnT7GPm4dv4xxBGbkv5qA
f4uz1Ko1TZYpHg6RonQmRj6bNaO8qeDD4JaEt8AIydEn2YoNHcxnq8zbBHjbfO28
pOiBn5O0S/7dxkpFKilHAWmw3NzgNnGEejcbdgzMEVX0wKoKna7muchKdouNua3D
A780UMeCSATKrQtgw8JreAmDeRaIkamyQsZHlAe0QVvZk+NF6FBXfa+U0z/URgYJ
7flqYoAzeAE6nUg7yKI4Xk0ljYhWh3+WHqXPK+V8kHKMdDkm0M4V0wYhc46KXGVg
DbeXt5kmleq2kUv4Wgk6Oj+6FQqEJuOwQv2cJyQqUo+aAqX8+nSFG1sE8clb+b5U
yxYe3wCFaVKV22E3L3rTDnEzKmuH+/X3cfW4gz+2jsYxMl/RSWxTPJ9UUxlITeqY
vXGjAVI5kCi9Ku9ZXDP1Rdbdu4DN9CCV+OwKq/a7HdhINUzsnxqNvy9JUeHECdyZ
/gDGccBeeu0xB5UCZm4WC+0yfcHUd+PNXXONTDBAO1PTldy6JfyrJI67ecIF8eUS
cvUf9Puksq7efVbWilTHI1d5xtNkv97jpYSojrS9fMhAL7STFW8MeELwTiLHZQzu
6AFGEPgmhjqT0mfP5PG8IA/swurMd3e9ezrWNP4OeLtFBievNGr5c6GPJnUTJ6Pw
l812duXIfQQP104mN+32lwmsMuW9+b0+Py+lB/TYlEMfgOUmoTRLP6PAmc61Bn+u
LUUjH45ByVYZlaXxZcNqMUDncMeZVh2c3lOdX3tWH9s03/CzweeWm2ITYtL1Maoj
W7lvhnuJPCdIBaeZLvLu5nkkXUid+YFextyUvXtEptdzTcL+9DJ4cl7grpQs+uoo
uG1l7AJuWSEftCcFTZpbVPRSm0WqH1ZM0Ej828ZoRHmNhRABVlaxLB6jyUGS2e06
Ikcv4Sw33EWrnfBIb8gc/TWgh+sDW20nkXRo6rBdtfEm7TXz5H/4k/87aMpZMwG9
1LTaCw3pb12Abt3puUJ+ziaZ/7GbXBhUNpO6XvW4+Vtbw0HtnX+uR88u9MEEUu6D
PjHM37hRvfA9NH0hUJVpryh/WYqtnudCgszAVRkD64IaI3XTp3HZ7rP5WcC5fqKm
wcJyUjxlMdk4T4OhlXYnKB07yIxaZraJhxt02Pdip0fQEv41f6otETN6+pGxLcQF
THr0ayLhl64sTu3xBQIHIjEUiER7j1KMjTl8I6RTQAecYxZ9CiM5mQLaYNmEhbNw
nXN1BcW6zWhg5KmvY9TxFPmUgLEgJcBJ/GMFHJ+pU5vvbDv8oJQhPvYfVEx42hT/
rpWRrokQkEoFU5qpLNwiQ3y3+cquB6yeMCtAXc1oqumuYrrwvy8bXiXG6GcshjyK
J2NXjzZM5mwjXQhJd+gH5kxzq6gwg3/6+3YUlxFQ8qbgUxqrgLBj6taljGs2U39S
qy+asZ8m6LWWpv15Dt2s0K9NF/4V7kPwxPCwX3G9nyQzxZl6k+W+3el/9uzE65zG
WpYA4OSaqRAmv3n1VZpeeGZOllf+K5pgnA1nutOOmT0SDbUHcg/Nvz3fUjfCRwxD
YpcqQaM8rX0VPuYhmgDkTZFycYmc/t+VdiFlkVWaQVD7Lg9rq/w8q9R6jsVLyJNQ
vC6r9G+0EvNq2PRJjAAJxOLIN7/MPE5Od0FseA4eidlMPD1SMywHE+Yg3BFHS77w
MSte8ZOgn5lQ/LJJyZpGL2XWdun/fPQnzSsv+YX2Qc7r3j40BqcTVJ7M/TDYHIrK
aWk11/E/iFWjCV1anYrb+NTDEPaHLvjYxh5fTuMtn03+DEcwpnnYIlYuCY9cI+M9
c5ZVBdKDAk+vuEAAvzm4xKPWauyrowVkJth6iTGpqHl6tvibH/F8BHLdwodViI4a
eLlXXSjL6lNhqPo6vutWKeKlUbKFDqZSg71Z3TNzFaAURhwDQwFaCZEhlu7eNK6D
sTtbzepBS4O1u2Fpenvyk1A/K0RTqgkB/b1JZFw81cCOZOcdPE2e1P5lBrBebo0M
z5XHYI9NPf0kW9xbcEK7zSasde1hr/Kp8Jt4bn3XnwEI0aWwJvknbTDh4QlrOpDB
9H+KUZko2vct8SqrMELUNJ37/3KH0XsiwQd6wO0X9VBfd2jLWBYqrXeMkxjO8p0f
CuZv9ehkJibzM4Vt91Qww5wSa5u6Y9pJrJHiLUamLPRKP0Umxd2qCe2qqBG7pehe
IviJUYeo02XiVFOmPBqYFVRKf+x+SfGu5XnLQ9nJ20UU4sSlB8TSLfj/up1wRQhI
dpat26/8lDVwXihxebxOKeBBGnHtjllU5E52zNS97mqs9nrkBLQuHsAZiHONUdk1
u2L0QlEsZbUH6ski4RSn7ifKHbhmZtpBp/OC03c60ltNMowDP9+GIaK1MVZ7y3Da
W9zFHqzL0TtDKtCRfj1neL9TGn8ojjsKbAJMDCYZaTdRd/OW5T9gjmpANztFsACr
Crj/tVAkBD6z3u969YMX3hljuv8jfGC7zFaUPJITv60PRcIJNAOr62Q67olSnA6E
4gg0NQce/RomsTvAtA4A5lGO/rMO/F+KWzBAiZ6w+TTAMYqwjVIHlYzpVVuJPi/S
jB4s4Sq7cdCw/Wtm1e8vEht8EfDw5Wc5YJPwrW8RivBLjBWvIpDV7IeFvzVl+4PW
LTDMwnVblP0AE9g0TZyC4tuJp7gr5sMkIrg4iIZa6zV796fFN6HxLJuOzih8cOb2
lG7ySedzUK2hKF23f0gjtBk897riCWSmsIzYgpLPjHRKm3KDgvsqSRk2vc0EqVAH
pY827cYXXrx8/QKhHIv3CnTg7m7q/Ane3OGYqBByCHefTug9O6v/z5dufUrnd5YZ
BRB/q1g0WQg5Dj0Zynwc2RHelF+snbAAxbmplRSUSHgb/VgVNqoRnDp+RrlL1c/e
3EIuzjkQMuDPmbz6X3ZcxLemD1M2mEMdFouumpT+KmIx7vitwoYe8SneeEy2yRVh
lC2rfC7zwJyDgGKemkLCZ484w/8kABWPY5ZRJ4OGycnSpH6iDqWWTPCtx2fRD+AK
L6eqmkSWq3vds9iNz8x1mHXZvPH1JWHd7nMLbGIsbKN/o9ZE6D9z8pam32Ya/NeQ
vPAaENu6v6kS8c0J41NH8/NqBIl+Pk2Pi2yESxxXUyMNuMR87KWuZxUyq4Zy5c8/
xhvTSJ5Wn4he1h7aH6gcLhuEbYK4e3rL/ZLmyOInyR6qSLrctayYTk6gylLz3kkq
v3XpEC5QbrvWrZK/jnx3aoskb+tGkUjFefKE4twSAQbcRFFrvQSqS3R01AUJLGjR
tCyxmOlNEvB6epyNJ0x58lWs7hqChZQstzP9IsIB32JtXCPYJTj4ynx1HYXK41Fv
D65ZPDxgVBC+4QWbZeH9j+m8NMSQCqmzaDxQMZRMUxNnk8NZuPn0n3tWtTsoMXxX
nZBGE9WJe4515znn25LbuObtZw81uUnQBKB85LSrORg16LBUTWYtsD1Yu87dhizm
8ZgVPCnP+o+OBEIwMHM9EzzsXIUSMDc3Se1YTJK23gx0/MqTaYbyqZOBKXAOuSyo
QTsdourHvpJuFeRpU/0MDlO546AJwAj2WFrDrji0QggbBV8zMHXwzhAGYilPZA4T
tyvHvTqxAxgTpSYfUOtrkOvLJq5DH/UgytTeQ//CzHj10CPg7wIn2B7XPdKQ+t6s
yNkL/J1UdfnVjSEmkgNHO1VNWijr9W3cZuk6AM9WY3Q096mkhhq+as9y1enIRzWV
TCvb7koHUWea11GFn/r68sMs+WAw812BSn2yeBYIbx+nLgVz9UVaWJfWC4Y4297V
VnaRwEccBa4rHQZWXybxNUsUFL7GKBeAcNMZe8yKqRnkL1GNnN8CXgZo1tEE9P9S
bQICHdgRjOc42cGmve41im5jRpaxy1g2MCfkLgG/YJtCCK+iHOZVOtb6jA9yojNO
o1xhmshHGmM3pFKSUMzAoEfXCUDcyhMiuWKBeVhhaNbmF3PnLVLSdadF19BhF4WY
Rb4meFJqSoYp6Ni0raCprOfzT1fg2gtNLYEXIOgVZ2g3ZGxfXCxrHb16pBP1kJwR
ym8mu1qalFIEwSyBnc7AE/yOftCGSWkyV2OE0EkA/VBG72xP20+4UOUZ3AKKUkCp
8TEW+IMsWmd3lq9FNPCrS5lUaVyTRyClrSSJBFn3Q8Zywgls5kJFcgcSVH/mL5+l
Sd7aZuiCMXwgb129AYuSLYB3rBpuCgzRG0upQpghPl29gSPvvWUw6zYK5+Ged3RY
Pnbvg88PDeHRmu8J94mvl3W5qtN01Buz3dor1d68LejpldP8B6I37NzJ+RPeJvwg
mnDAwVBTeXhogf2FRETyzfhJuyBvmGnTxwN+w2lnNjslvtQnuFI1X6QqVky0syqV
ln/ReCSmvKNekvh1xhDYTUXsERJdwrcs8mHJMHEbzO66PIy7UpLxnoK0H/6cu02F
EmSJ1fMgHP6qEBvgeQsPrvsWDtIPI8F3iSVkbuVSJW0XTY5N/zHmbzJbjyGQbbGr
pjJXY1ft4t6uDiy2S/rkqt91xWQjStQMZrWytbb+GUhGD8szSL2hikKoCWyz/JRj
m9ClRKlBpjvW/foRLvNij++SpeFKnKDyR1HNrV2PSRYWoOwmDScJ+nSEovbb6ztu
3xAGEwfbfhxJCEwprml61Gmqpq/SH92vRIQBtVCN4j9+KbjoQCncnbVE/scA6TpJ
Yq4su+C9DUn1PU29+wfcrLkrSSxwHRzEl83v/IR/rc06z7Uw0Gq5FABmsfKIS5KU
vYOpFegX8yETZeW/rAQpMO5GKCY/Y06o6MpCICFk7SIrugUs8dQ7EpCV9dj6fkPi
rYNRKjHJyDX+4qDNG+4LGObNO/2+6OcjuCP+VGdTsXuorQt3k0D4p4Tfz+x/c8gD
i+8RpVXdZTFkqx7bCiRQlwkkVDCr23tU6p/Uzej+/6lY+ZV78ef2s4xcBt2Fj0bW
ZYdRGN2aEzGTezuEifFiCxC4kMQAL2i6f1fYIr7zNm6NFiT5LkyhhXVjb2TaLd2s
RENgZiapi5P1lrY5zyJGT2/Smp3aO4pNuLrLA7xckn/O//MiMJX4aIjQBE6ZvTfE
Yr2OnJ8zobJUvo5997saG+EvpMZ3vpHvDU8OrGAVujRERcHYUGlgEaeHcd9orCsD
zgRUcMLjQlooSI1P1DWCezH8MAT5yfGZPqfRIclP0iFqTvEAbzZdvFopDQ5vvYIg
6uccQ7CbzGDonjpWWOnb3TpobaEk++zZ9OmGp+X6VnUHtqJs4JCK3hn7Z6WPTWke
bm4zYRBOkYZZianRNeClMPSBk3jA620SiZTRanhfuY/d4Vo+5//7XI5xotkR5rvI
ubEtV5FfyllgDotMNoRSXGHIm9sVUd68VJBJX2VMZFjjrByBSjKM1ImsHxXuoDq7
MpcSaWZAH+d4gZNO7f9uBw6Jv9lCs7c3VMZ17fA6VptWJ7T8P/rK06PolP+Y+Zvs
VL3HgKlhcrMIrLVMlggpR1ebACyb2ONZn5TS1VwWRZNlQZ5C75TOpaGQhkFbX7Ix
hQCsHQAGEN5nvEP8+5UMdhmQm+pAUFu6D8wIVE5VR9Hq+mHDgC6yGPgF3IhlX0t6
dNvcTVOHt2vE7vZpCjNL/Axe+Sll06iC/YUi+is+t8Q/h4H0FCJ4Fk+xU2+HXsd3
LbzGuLPZNKx8WXVsy7jlgLhtsRTFvg67/AHvz9nQepbtZQt8Qu2AfUWsxn1DY+qp
Sny8ng3EwzhSMIIMR+L13ym1t/MB14FUm1ZQaQED3I9NKWZNOU2BSwdZUlfnRctC
NoMEmmD2CtfTDN5GIdv6I4PGfQW42wgCB6CUtq+IUN9VoE4E6SjQTozTYOGyCc+X
tv4OWYQB/bPqP2uFDeOSB0XNvf6YysiPqRjUxXTQAPSHXuwKqHou6OdH24RNfkvW
lUaVquMZpT1SmNqYMW7jyZl+jvsU/koVVkrd9iQYDcJHBsFmCNO0+3p1Uwsb3idI
jNYnOM0VGAtr5WFMGcuJXMYLMW5VW7UB//5LKzePkUNVsGbuXv2KQ5mOYRSzTUqL
KTcQM4qpOSSdM2CIioytb8lq2fuSXsRcNGQt3EDtayAxi1QNcoOIQotmyIBUgCFI
c+/hhezjn+Pwuraotehrs9+fyXoSuVvkvw+E9H/lkKFXuEEvgQmfIbBZNgbCFgXQ
BKKdB+OA2wd+frSgj/3Cke+q9KMkT//+iurA0K03FAiMwSaZe3h0SJKO8oICiyOs
8fOIEYHX05x4dI7P07nhz/S5DXYpZra+Kpt3YnWyDmZ+M3MEEWBoOoSGySOmKSN/
/2QYFFKllg6HclI7Izs4DO6MpRF87tlMg4r2D+9yeyANKLS+ZGXEdIi5t571YyU1
cIdkqKDlrolub+5VieouqaKFkWKFSNeBCbPo6vz1HL4eGDDCUSTCn6O20z3EgVrZ
tMwAqGYYkKV4obPf5BUx/of0bSoKa9yvTJY6rez9ypxX5zTNG20b+fxp6A81DBh4
icVFLXGdOg6kFTTXOaPtdhiuEjME5MtvJ1IhBn3J3D4ASQXVlsO+ceSJUEyjGVYH
MGmcb6K57oHaGFKZHkmENyorliIoY/j+IeB7mwNo3h7ONgBVCHpNYeT1gmp23Mj7
GJFv6C9xPxZZrReUMp8PB6XSgYsuo+pdtYzEt8n0OXhn6VasPH/TaFz60upujnr/
Nx+Fi6dnpjpfbA/AFk6mHl/tn0pF/2Z16qwpTeZiI3D3CkedaHY73jBqoYBmiYsQ
IM/nfum23BVuNtQf5LaYVnTRoMY3gelgJ3fFcVRIM7LJ6nEnKCh2yo7xy/EsFsZX
jzuZkR8yTsOLVncJH6NFMGutKLo63LC9ip2yASRVNlYLiXgjc1s11qGVqnTi7d1U
fZrl5t7hMKdzMhAJsy0rkzt9G10+pTZEjK+QZX67l/O2kAJNdsaTWHIMQdO+2XwB
Ax4XN+onnz8mqQjiHd7jpwMG1f4Kij6fek7afv6Tk1S162ohwCRc1Z1wnJuGB/4K
CwkBe4WZXEBoANhQjsL8OTo4gzK8vwuDc8zgqXYjYvFlXInPerC4LviZO/Jf+D8v
sTVLXrvFhiMzCKpt9Dbv6LanGSULyPugs+55rbZLcZSJH+uv0DnHEXUShHMZmVVQ
+DMOm7V6vjyjpLtWWVtAM4ud6RevKmgg2HDZQaTjQiU453IgGrJY0TMo0lQylUev
bbEETgOAxgUcQll9jST+KfhMISTdYmNnJPnFryZlQAbHXTSqL7wRHmGPW1MsQvuJ
HjCBTLQ1GVh/2v+R11CdNL0KQEPEaxyy6BhU5n1znGWRMYh8OVNS6noUX+0lXR6U
ND8B1UJzscUCK/IoBdweDpfKZttj8a0FJ0ZMyb3eaZQJfsl1gdS81eHIKkB/4u6J
aeqw6C/PKGIGOd5dRTULwrJ66wFUbikznxY/IaD+fb+C1j+xIlIT2ksW2muGxFXM
N1qAOqFrAMbwi4ZACXo9Vd0vIo3E+voUqHdI2jS3b9Nt7DiAgGEQsZtiArdvEG9R
lPiuc6+apq0LfEVogkDYRJIxU1Aintv6aNsbYdFYx8QF6c2YrJJ1IqSiPr9pI9pn
gJAl/WBG7Xr7GTZ2/m1A//wHKE0N/52R5TzqdSxwBm+2KB46Xuq+8n7HUDioCjPH
WoPMwu+HYAQWEZ9Ihnwfl9+ZLlPia88VEDD6Z+Lo8juMG8pWtZxBDY6PO4eGaWuO
tRga+RFYVGCnPn7Yyb22sm4kfk35DpWOYMBWHyuNE0Yr/uwKpDzut59GlTFIvHvE
r3ndI7feyw5jQpRNzT/9GLW37wl8s+DvSH7kHglzX2XeAJF2JykmivGFIJS4nTLI
VTmGHpTlgOLIEs/n5aAFBdSIO6QZY0cgZJt71l8p3ApBnNKM2d2k6ICJ8AAzZJda
jB6BvBkZ5u4xQGb1LU2aP8Dwid8WeNMgDgGzXe5mRww6HLiRFQEbAsLH23k7a5d7
VzKd243j2Qbl9eyA6k/VQYqBEKPoThDp/UqxNKVaOblvmckLS5ndxMy/ju2ut6ZJ
JJ9y6aHRTmKUo6J9DKV03Dm5+moFcHF0bSOXJ+KT4vAE62KhasLjRy4awePwlDxC
Gplh0Bwz6dpNB/rx3rPV70DcaUVbxbple7VpC/O2MHmSemTq/Py1fuWQd+chpZsT
ms2SkmKBOn4QgRurEVA4zoi9p4Xi3sjrWp8KsZRcXGDNvDWo4COwp2qB7fZUNeI+
6qTSgQdI0hswIc1EpVe/NiJfDj5FI4OnbdHhhF2hUFvnP9Uj6VTOOIwSK8L0KPrO
CNrwX2hq96if+sEDMozdrMG99XWw0N2Kek+B0XEiywPayvZ4xeF4PzvBg3XiJpn/
Ew3PJ/h2DofiaSH//9w8MuMMZXzIS3J15v/h2FMnDKJFpetC7uvbrYoCEAq8W/m2
/m76FD1vVBBCxOhpsc0PQT4Yl4P/3ijxvDhtF+mxvk6fNBXbPzdlb+ZVE27chazo
/Jnzvdrb//hDWzRN/3xoici84h9ceGJNYNQpMNWcNSj5htbEIJmAcl/u3MPETkhW
D0V5De8uBEOwrh7JD+PC8xLJsRpnS21Jh09uQqxNzTM3ptL3+RszfaNes+7LI5DC
oo5AMbpnZWMqxyB2u1c0yotiW2qbcGze3M9fJR2E59A/CL5Ec2A92vdYjzyYe1E1
PXb9ZssQcysJ0FFYmaE5LmcVMrghqG5usYrZyiW9TomiKXM2oQH1RDaaPgiGawIQ
r8a/pGsRWokbSkvs1yudEbUjhwNH69WsWC9JnWrhVroCdtvw2CXw+NEjBnoRYPgd
BkIwgJeG67/chfzCDI4X3FG4Vx2R5I2YgcSuXQQT7BL/IULLTFuiE/OG4kMC5vMF
C1JOHSXJfbQhVUBR9C1bGZY9o1u2MGsQgDbdkKBpIXN0zA0S9G4/6nLzl4MrbjD/
iMgdoDOnsm68lV1G9h5Bw+1Mhtk3bgye60xpVs1vFgOFh3boF7cpNaecZ2lyyAXQ
QIjKBJIT5qRM8jcCkZH7tnHRV7Wtw0UTM4/eEHlSpv7f9Ug6uUtCYbEJhGA4O8rW
Wd/j0FTlGRinEl2Jxcpy9fhmvxbWYlqUzBH+dGMKdRAu25cE7m92HeC6FjJHMhIN
rlVcB/zdhVmtRgN9jtwJxqR87WUzyrLJ8RrjQKTH8oRZt18w+1L2zRcFRToG4PTV
9/Dx2LLs7f+HdQjpvoRgWH3wxhdw3+pZwunoJ4GcHBgC2dnS7HHWajWoHHGUbRjy
rpAO8wq3IK+gYvF82+RZWKzkTqatM+uzjRSdBNYjHqNO91QbDLUyyvxfXk255t42
xT0nIRNRkAX7ntdIrXQSIkEK+aS8zKV2MBUZJ9r7kXC41WjBIdi9cFH1jw4yfGy0
mz9/0VfRq+KUSKwmUSVyLHEKvkMdtmM+Y9aUjGTsZCVljtYm0cffqw6A0CWkbDJt
SA0dtEANQV4cyU7mQO5mIKfUfPEvz9f0PvH3pZKf7iVBeH7pMUUtTL4975qQq3T8
TGaDnafgEAKojTYvSQ2KSyREbnb+K2n8JNAbVdG2pbVLZTZK1ZAP0W+2Sw+laFxf
N308mnqzD9EWViRDB0ykKelc7lg4nVBMLTg3C6iGs9ykwTLneIjJgRLl3pSpPLeG
cZDCVvBHs99mGoZk5DfJ5myLEewBdTPu58w9Tzns5/1uxFR6jC7uXHUfGhZTHjyE
EcibEi1FVkLuc6tL888klhw//cZoCzmpS2w5ADriwqjpk9XuwwIdWAqlGSHnsMff
2eDnv9nTMkBGhIEk8ERtXI7ow+K0EE2SezHajNCnv6JQf8I51tiHOLaCMrgPL57w
09Si0IEWUmT7JwzRQEpR72E6C2PIpx0Fco7D2bF5+yQfLTPCDrFnrSVRLdYurkzj
4W4b+mjsNio4wMXULDHvXsGlnYwbn15Vqeb6zMoumS4VwhhXmR6+38KDItjyQkC6
Ryf0G/gTYNSHJSi2pr2OEl+p7ECwU3KBk4DMDJA1yb+GVMRgyxvWU8R0dnpLNgFd
MhBqRGOTaQ1lDerRmWW3xLUrdGLL3Na3D24ubrlSrvYnkCXE1F4EU0xWxwV5LR31
6+gwzEuai90NdZtrfp4lqHwXflnNHBSbqYmdN9ZEL+sfbwgrW0qhPRw74wn9eO4e
wR5uV/21Hn8kIWwCtHlbWPCKO95sUffpW9WhAdidVV3Rr3AjXmv/tH50Bs3xngNR
6m4LZwTE9j72jecTMcUhoAjHqe6/Wt0JFcZyMa72fOhn/K3FfpxDFb1nBMDDFf2A
GA30nZ8GQtKtkXnApAPfW5AePEzcCIuZ/DlULWAAZ/ZjnOVSaQN7EUIvjrVAafIE
vJOfsjAipQtCtUKopshkChwfCS5SMcsMp4Qp+Ws0I6cAy+t/hjm1ffvEO3BjtPwm
Px5KDIeUg8mLlTeqcW1qgIant+M5aZ3LwJoklooRTJVEV4fZ9ySZrAW0+YzaMSZQ
Y79GAeGimWOyCYalFJo+t38n7enwH+el6sE3sPxaV68VntqsUTGK5b0suL35guGX
d8WRsy3uWYeVFRz2PcVIzu5/mR15zM45jfasaEsKSX3Bc1w0FGtrhw3sBkzq1SPz
ojdlaPc04k4/d4KjHTWuIuhS+xdMurtTJYiPAwbyczMOvYdzis7dQnYn7RlCMtgA
H3AIRg0zEpcRcLbKNXY7GJbRpsOtBEJrxhuf56tptgg6M+jge4CWztOUYQsTcO+7
ZV+INL4+7C7yFe+JPWxrRujSK8uGrji3YCikpKIJTDtgh27QrgzoZRKsBXxeMITF
ixdLCCgtJsjV9mDjwv+M++820zczcRn1qOUlRpjsr3o7LRwcnZSXS819OsDfMEj3
sZmVUUcOKUFqxzAdHEd3ii+tDVKaG0O84FLREB68IsVkJWT5EHE7GUFt0zPBjaSk
wA0nNHGBJwKM57qrPtAePKTnv61/waeEkQO6eKXqrZMkBwER8x3PqG7r6s9SQ3io
G71wdG2jcgm5hEBsLpywiLK5m49c1/2qlguDPcQZh+3nA88P5nlvkzpwZKV9er9D
qkTS4vRicO9WJkinuxYyItF80F6vawY6ATL3/tlLOfVdjGbH62fMWu/IpvVOrwZ9
0PYQzwqUNIbzQSvdfy9Dh0W6VCRd1oa27es0u4XesHGgW6MODBqXhDorlhs15jQU
SQbtd8w96QYESfZCYR7Q82mFPtTl7mLM7dnKg+jQCBncetU8rlzCjxhUeWTri2K0
LL5IFEXVOG7QhWWL8/t7cew35JxTgANEQt1Hjpc8IJKTWiOkcKg1mAs+41yTDeHh
6eht8XEvvOiQXXiujaAZv9RnE5UKYIrAQrotnndx8Z6aEr3XI2GAWjfquc8rX1Lm
wZmtilLGWxwkzShq4sliY48OjK58zPhV3kOO2hrH+j3ihYenX5Y0vpxlSYoN8Jz6
7bcPGnnHuJi009XDagmjEdCL5hQBkcma5FHLZCdYm4b1/fZzzWTdJ/XO4PayaZ6A
lPNz4UzGiVk2nfBT5pTbOw5CWcfttYjwIjBhWkDngkyjxUpXi9woE9MKu6d71Q7a
xvosF10aGaxDQFXjfShGmqq2SZ59hgeL3DhGf1Diq927UO9lQDLbZeVK8BFo7eqQ
VMecccmrt6fGZIFpZMPUYTAgDUdzfSg+jdNOzXAOICZx/olOYKPeZHP0qNRIaNSU
GPM5bZuDHjWU58vRjehuVk3tUrR8eYYEEbKjstSe6stb0yx0YztZk6H05ANLYJSC
Jjm7hNMjAGR1hDqWjdFO0A2SXBpDgl7yaaWm1zgeGnXQnd6mgMFqnBlS6E1UI5FB
n252f0AwXwTZMJ/y7CC7aRoHXijjAzZA1D/3oB21QaEj8Euj2nOiBroT9JfDbk0y
Tg+g0Be3XZhztvI0MX0PqfNaeC2SQiC63ebF5l0y9/8qpVHqibUpUOOZ0j1gqyLY
+FuCzSrkOd7z0uUj8cbcEuCedwY5vZJyHOEkhMn2TDxWgKWTNq7soqU5dqFKAfmo
IsPrgDSKHSddRaOoGS6WiohZVVdRQIHZeywLoRJmm/c/yRjy1O8LCVRxOT5zGiN+
UudHb+fy/YdwI/slqlKQOyIA64/FzPsxn4XCcEIv1FugLT1Com6GX57ypbePfmhk
08eafHo2IZlfrb8dzNNu1dDr/XDTN4/BmDpIsJBe81Xq1Ue4p07pcqu7GxKeBGBb
B2a+mFN6zM2+dvgZ0Xsr8xEKEaTu3mpf9L3cQyeAKb1mONr5PCBPsP6jqoB1yR9K
Am+po88QBGp0dOfnO9+Zdu1opfuqYrZhuUGWFBRtS6RzzRSV6QlPTVXij04UU/dG
G/5pj1nn0V1Xif0joMhxHdudkACI0Z445+zLH+EnZpoePdqc2bNcLmz4cEgIKQdK
5Mr2o2bQY7Ir/i/glAm3BYdFI7WnyFJJk4G8SuWN6Fo/zEY/aRt0xZbW4B7RFNit
L65RuoJ8Ekbq84bafvUMmd8H+rJPsZ9AzDvfxlAPms2GjTNRTDkeOGkOY2bXtxn5
ib6kkKYHk+dtyf81rtmtVW5aKAmKEduePjhCA7eWIMQ30jwqa+jXhksRmol0nVnB
ezbRSgPSkf7fuwhvgY3jj6yCtqXnNSAp7JjY1X3qqFwLlQabsrWOW4EnP6PEMaAb
VOTPhC2jAsSj2OgQQOn8ZIsEej+GAWph/I0ay1xw3heo+uYKADMTiNktM1zS0mTI
4+VkLhI1Wiz5ozUfQ0nkKGFO/oWd80/YfORuLhgU/WdKEy/0toYpOgl3yTGH9jta
d3RYaOOGz2wGYRlErZ3Rb2O7o8lq+TBMqor6o17z2utQ9iKWW7H2NLxxksGSB5bG
8J0RFMzrr09Q71a1l4Rw1mHeU8DqocTFnbZP0904cHcwJIPFeknie8u5C42w4kPE
YAaPHFajarE+jkdId1ZR/EIpQsqeCUd7LoPAAPC8DLm60dGIOywGRS/r7d0UVQDN
8MYV4nWzg7rFi28yg2o6OrxeO2/mETDR2MGR+6M2e1D1RPBKg0/QCU1S4qnkjH/g
AjkY6rGnY99TATBB11DKzhEDfEdZj35rVYsyzb+fjFCxJ3Uv/WBpzEOGOnjJ6iKu
CbdnrbkU5Z52xYY6SxuEYRpjuPRbTKL7tQzTyQ6OQIylPMEs1N2vwTg+Q34RhZk0
2sMrZuch6mydw9b7VEIaEeQfn/2O8uwZfy4DQqz09a0stxFw4XIQPhuBg6d+8zru
Y+OAfLd+ciWPSxd7JHoBBpwgnZ0R96yH0D8YYdRQcRy/IYMUzSTusAa+3ELY8MDm
f/5yZRj2Kcw44W69z4iOlJAnNQrJ9wVDyxJ71aC65suWpO2RAqblorBA1X/5qpkj
9rye1oI3yWliRYVspwKPtx0x4zSZqcGvTbBRfmKot+KNdujGiSUbXGUY9t/Pkj3X
SdwejjHtWskQNZrgjkw2qKmBNOWu3N9xjZ1jW0LU/riWH/CJlDCkdzl+5eZTmuaS
3I+7d+DP3u0CudL5ByYfgPPTTSuHMP1J4nlJzoMFKjJdPIgWcVHaAxtZtKT8y4w+
+RYvaHDeoYc9gK1gDnClzKBw+7CT7QMZTQMCog2ld1sr8CyaOTUlQTa83U7d8tAj
IGTSl1rjBRm7l//U5Qi/clh8SNUCCgNe4br8EDkkuO1H8SQRtjBQ+OFyTTRLhjw5
qdMWCtIRbz5PS20tawdW09eLo5mN5sVaeFHtfsiDwez90dH7xUYUumStE2sunrKL
RlmwbWEpMl10T7mQwGY7QI8iu2adhfgOsw+xeGAfsDtwseeb0XIAoNh1DOUTlY8F
DkkbXVq66AmLFVWmIzKOxTbZ3KoTF9Y2YpmuPqmai4cVN7mIheCxxiVCHkYUYjRC
TeuRlKtADECKszV++OYbYik2tj1T37LcBTTYo2Vo5wSVgMGL97UfF8lNTZWb5fYe
kbdYWG4nGwhlWGnYSRmCuKFtBhitHIxv2KXrvQLWy4yjIReSN/aUyYbmg4S2PLeD
Va/jltcSC63bqQgO5jluTqKLscbVZ1XImmFFlWxSTLBvLJ14QzTquKOXx/iqIhQn
SNgsFNRPYj5+Rf9F5sBeLG1iY+PxhMLNwUYYbQy5KxOjpUz6ceX7CeEYnVhtcvdS
pnzSu6+Ltd31fSy4bVFrdFOmVqSGIcu6OMgvHK1Zjdjlf1l2JiqaPsgcV4LTfbHF
DhVOg6pkrCbuRzJJCh3vmtQoSnGDkoQuwrjzNoq4ag5VFyXXkRc7bhFGS/b/BD3d
lcxWUhUEXHCvEG1z1VAnEa8x2OjigqEKk0s8uBwSm6APO9KU3X8dsz0f6wGb+3gL
BcHvkMnUHn7dn8xPorODf0Z0DqqJ+veEdhYZ6Zp8QCfmh0TO4kgTBNPDcIvDf+bL
AoL+c4ZLaer+j1+dK5AfaB0Ao8BHLloP/8YQFX0wtGGwXsUMRUOwxGOmm149biay
WyjB9xXeMEVWNI/XxA18Pk6n0m0uXZmG1RDJS5s5DleIuuPpyyJSSxXVWJd9nb/q
RiKDRJenP7HkhKv7JV0wym8x4mHodP43MiRjsVbkSFN+XrXwaWo92vcrF1Gnu0M3
X/h6vyU4IEQSfe32OEDWt6rppNfG/uNbZQpTYjVz32ObUmIz9vN2vr7AyT3RARlO
8E5cjus4cL6SQrTB7YY17Zur2WLJ5a75LuuG0NJTEDzAZa8c6EubiHtOfAnASC6/
bifCtyTTvUcEPJchUoEHPiprWvgFw+EYvaAKuhSsNXaR98R2bZqjYOJ2dAoREZHT
zd/wXvX1RykBfVKq549i34rpF9qNEPXtuzE0/lrdSUmEFwN34YhWTq856mxdLTKY
F6EAaNGNgLBaQuuMTw74nq75Wn0cOS83emGGXY0Hw0tKxhE/WlofH78Kqx1aZgxM
97DZWeyvZgJQRRnXNFB3qMEWWo/sOsp2F7LByjc9FHW0kpL43/KisVZ+qHbECYXb
6zuqYg+5avX2B8BQ10nbQgC6qtCo9Yl9WXiwSkAtG+KeFvcmyX4rK0NNsXRVEml0
v2G8EYWVSuRompvw3dUm7ZzZBns/h7X9MA0693erVBllzFsPX3ZIsUajrzHOWYEW
e9RfdW+E9HIaH6vuRl44gyYxml8+n/gZyE/dBR4J6U/RVxe20bTKu/IQHK9tem7V
6jGwR5Ju6W23J4uu9hKAJDqiKBf4mAOIGA1oNrfMiT1slL/bm4LxueF7ZsTX/xfe
ALyfOzfSljMt+s0BECbR+pjGIOzT/14xkdNimZt0vOm1yjGLJ+C1mK0DPSYJDOKA
mNKOWptnqfrMcXEa5f4THZD/JGOPJyq7+djXEOGTv3fhaXsVdl5xZ3dkdiS9o64J
qNbN+qxjCWFzIIj5drx/SIabOXX17mKYsCWB33/KN+2KcJnEiOnLaQ1CS4UDRMRT
beHIo0LEQeaRYDLW50wjkI5SITLKv3ux46rBtfetJB9o1+28r8K9LbX/uHAnaiX/
eKwgRk5qNNiW/JD1O3nfO+luTisEdZhm58vxsgDKCgEq/XCFuyAULo+O1WFUDUCT
zl0VkS+hWzOzjZ2LspgrkwoKJlX7Bwhowq5eFckRQTienLvovyoT9oBrpd7d7N3S
NoQwGW+LK1SEtKV/WB7pm5nfl32dfwFCo+UqpplSAtXXaDpHc1aP+3GQCR9Kwje7
ZHtgNWcUzpC/OM9FRkwOs52h0ds0fHh5lUqChXkCWTPzwMXdXJ7+gFPD07f1QUpe
9Stt3sh2jZPndJBjqEzPQr4zpkOANXUklxqKHDNS2KJMY2K7BJfUZDs5HhGpS/Yo
1yYz5mw9DRql+MfUiSPMjL++AnhKoB7SzMf58yiTV9ONP5GfRzuT5OIbnvRUaKTr
1juXuSHsDQmoDcLu/4RQqxpj72R2+lESmyJ1uahNB532kT2s9OSAOHbewrTx+8Ic
LDIFTSDvHfNmkQ0s/Md6afCttgwdPmUKMWwiU0AYiN8S3YKNafq86EahvpfqLhAY
K/F4WlHLgKonVWWaGutC79sBpPO2d0nvkB+fARy1OJ0+QLsphJlauTi8SCmpmZS3
nrfs5QjLBQYdz7PMkwHNGKSqLRy2xFtP8xpY5I1NLl+m2tvU8Z51PCUucRk4NJTV
Zcn0pFj3jfkGRbkGoX4GxzvfoQypgH9Cf0/JiifKh6hVD74vu9GG44Y9hmTXMfZx
4K34ESnjy86JY5uSzD/VgPwqxRAhAkudNPuE4XNXe8IVkihx9+pReUzOslMB5sj2
pZtHQHHt2ao+P++6IONYcbWE3OavEoG9km/eXas6Zoe4V/4Kp6FJXHXYklKVT4XX
1VFj6yoO4vF3jyh1ZLN2iiijA+F9w9d3gyGCrTuJpn4+pG1C87YL5lzk8wZi7uy7
oGgmIc/5Dk1lY7iWaY/T2h0c9Lb4u3qWE+JCqI1rz3apoZ0u5NT14F5xF9dqvEsR
L6a3NL8wJCxB/B0aUJkrGG+retFMBS7E1G35YypyG8pnLP/ML9M/aMFiJdrWToqf
NHtbNYpY7fSBHUZTgQgIhFNmkoClhZsC8HYcQ4+wn81zsWPJ1ULmvECJsQYpt8F8
1tBy0diKCKJZEdto1ozqfnwam7lVzZEC95Iz/s569UEoLww2kSP1ys9K0ZnJqz9+
ItWUH0DZtPjr/pJ2czFUViTi3XZe8U0HNWNTkTgS43yPS27VXHyupXnqMQs2f8W+
4HlFMgh75CJsR5qYDH0e2fL+hZWiZbMnw+k5PMYwjTTIhNLT/G6DwxvFJK5PAhHN
i5biJA277osgtnLST6pdtCsE+yELw0FkZq/EYYU0xLiDAbDVBCGQYeIvgeXno452
ZTmICFl6lbxjPz2HXSHEYI6MEBzbuXHtMtIm6Vkj5/roQh/Vd70ATuyYjIpJz8NH
9ZknUejcM+vY8oHa1xziA7Un88LbpwWdFC+jrkjWeIhNdce6v4Mj8Qs0hsaNqioV
Lx9WUkys1hByRbsISAlWSyMbBLY95NaIdyLNXiTV60zNsmiiC0OsQLHgQpQ0gXAe
pM6nMQo5DXfUDYCFad0b23o07leSRR04kaYynvM4t5JkE7EjDRVS0wIXNOipPFsi
IWAgn6wcvKCczCXyX2+LyVjD/JCgcQdLNZQAyj8+PKV59G/bg0UfubGia4F5GDVf
MCEqPabDjqWic01en6gWRxk8tbT8lsWm2tFU+b5fxb2lk6bSIW4LuiLDU3/wTFYx
dmCEbP6feiHVTuQNkcmVHZfbDcE0lZ7Tm+lDICud3hsTQ1K3D93PsttE5GmzqroD
kF58Dw7d66CqzgX0ryzz8yzt/FwacTmMp7px7Wu+dURSFf8WPAyOcf7QVxE6KeYj
PqzT/tNZOOHuZuH9MaJkcp0BsWt6AzPfLoS2c/lAF2oJl/gWAReevxiLCXYI6Fun
HrrIgE3VxKHrHCONbltY82EyzbiqOcbSrOzlp7+EQ/RukTdFYcQq6lUM/ZJrEHy6
enaq83S+XDjlhtklTRCa5dufR5xDpoThr5b3R62x6vnSNAeeNxiW6KRQvJxh4vpS
bR3KtGn/DsH0qpazGhml2mPuVp6kxEbwuKViLNVmYvJrsdtpsPkDWOHJW/v0eltx
VWntrOAlrT4X+MiXJ1anNLoH3yLAPwOKtYtRq7XxxEG9BxxLvAuFmW1oro+a/F/d
HSgYv4vkmcQVBDi6wQziWggEaMo0YZvc41Ev48fxeeo0gf5UcVU5lF6Un2wDilXU
W3/f6gdXOqE1dDWZleb002btV+W/zq3OEp6kWMWA4Lyr42p4srFoEZwX0tHTL23U
mxAeNccdLzLqNMPcjO8cUEWufb8dL10u+XoTvzcJlQmg2BcSGRv2+5beXs9GX+0j
DqRu3VetHVQlUefwaQZVQjwKGObFcPIszSe4BTAulIcITVqNjIlrClMbC6SKUGw5
LM+Aa+rbKDcYze2C3D22deywIrJcLaW8sJiqAvo12dqCS8OuCSDbqPDXb1xmm6X7
HOx9UqWliokdGGUTKWbhlCSFbUe6QOicvG9WSM1LXMtD6qDXYoxjPoj4fjGPDeeU
txh1Bgv/xqjCJfaF1Sz0R3zcLBetNTW1vegZfYBFWbEbJKviBBCxXcDp2bZIJ7be
GIUDnWRTdz9DA+cfVNtKCDx+CHA3Mp9UCEKpxyMvo7XsFxUy5852MPr1Is/qe4pN
Hbh3vdlQ4LgMNBP03NdF8OT634VnGaHaJOMJWidnAAJsZIkS2Gl5QZ0hTUPxwk7U
3D2o08uPHHXvONCBLjGUuVGqExhg9NiPfVTjcCDegjyzgR9dfwWJiDrwc5rsXfMn
HhnRNR7O9p22RDSmfEtuu9dvq7Vb8LSlhQjJWxoaxOwFsAdvLorPDqF9SbRwJZtI
9i2r9+YxSJwg6CZz3s74bI29yQJeoyyHUg3vykoRQfx0/wSRi0Z7dkhqct99t9mN
x37cjKQnoyPaWLI8gfGlaPOZt22NqgE85iJI1lgu9e3zGma8mzuMW1gti1DOwhiW
kgVoPSbczzFX32MZOKKcD6br0sfwMQgU1ThJTwNa3HSi603piuINEJi+4a3TW1Mp
TNvTTBIlz6kG1HmS/XmDxUhomvsA7IPlchFr5eqVqrK15zbaPhzSjARTd8gg62ZJ
7Zak+ktaZY1a++rnFFWULzxfwbJ41QPP4rjAo/LlkbTdwOKGFRGKKAK8BUhm5745
s4FBsXPxMJQRp6GjhRjizx81ayWOi4SWVtK8FhCc3R9qyrcK/+va+je2n7PaTbmK
KPYken9DZQ8nvT97We5yZIeskkwJCwJMwiJEpoLICmtPNT0EcqiSYW5e5M16GTyR
iJq4hH1yWp0/+Ej6mXfmlcoa6gr00DncPWDPCPW3T7pEGwcWYOruaCY5ggHS0iys
hEmqS0WvgVVFg8pbgoRQA/VAKRfAVwVpLsH+O+XHo8b8WhCMm+J0aMsoJCTq5cBl
eWsttccZlJzWW5kqh3O24oAGCpEVRfSBcFgr/DDP1Pc9HfKxUBgbntLlCB3VMCI7
dSA1p6ydpvzv7DEqIPvdP8iNLFhTp2p84EO27Nf9GUvMftso6tlRvy2kfVWh9KQv
41eI/x2l2Ur/uK9dMrSIO4EHlYKG8FGtlg3/PtK44h4lW4DWBelmK82ve+lqC63U
LxlSET1Qd1lf0uGUCQo9sC3lUuIjR68lK9v68BgjcowYfvAkY3my2xS1y2eCg/pZ
rXfl4IjlRVRJruvA0/un9+hF/gY66vBeFCOMjB8AnCvZqpQM815Eal5ptIbMUQ02
eZXKpkiecbqzg28oV1Q1bN+g/gd4q/dXadOgE5GYLXaxOhQOLeDTABh0somwfwX9
CJWAVXIL/hDYWJ+9olmeF61dcpbxmhx0XrMQmRKDDb67rOA19aTo7n2fDiTOXq8h
plDoEMj013Lza+G3CF9/NyzHq+8wtmc3MYh6rc9qF0isuW56YS7DFjUjpHxzl7l5
FOMhBMvGgQ/jFjMGppitbLOD/oDbDDebyyIzVddPWAZPlfvSpbsXoZlsJZV9kh64
SUBeW8m7X4vTsdhXzrR0+iBrpvRACbakWhlmS+1enIlj/HOsnjaNrP4GsGljeEUV
dbYhFtM0I7JT47L24UQje3VpAFuQhuKLpbNYZyLx3MdMofLlqGKntUF0k9xLbZ73
Af9Zgf6WG8YDgTNBtMDGBpJok5Xr648BfQrxcv0Bc32bnYYDPibFvJ837fxhQMQW
JEMRuS7G6Wx8kVRemV7TwIhp6bw7WT8LnvP3opRlsw31FpDrZawKLFHyYQyL596A
8JsyM+ssLoP94xrtWXkrlvFH7EWmQGHD8bwRXGG0gVSTwB5QFupyj6GkaqzdnSr0
UYS0y72cY/7AIlfGVc5bJ9Ylz5v6742n1HejbjJpAdKy5obRmgQAEW1IXa5qfYuY
U7N1gF8ZjhntLc9dmdeufE2z/qcwu3gLsiqZQC6kMVi/pKVYgSaPM4zcsssTj6WE
QsV2uy+oAfsPbUZl7UzRl8OSCMaM3eRNGvSkp0qZMgpddza6XxTm88IUA66TKdW9
tHb/HuYdtnvBkmtH4lP6nY9gNZ1UxIRT8gaXhJ0bQQWDFMjUsm2DHwj/pu3Hkx20
yuI0isZPDQznMTkiyrGiK1NTwdw3jeyq21uC1UtOCbJe+ibDStW21r3kpOHsOy4A
dUWISD2E6fjEuOKo2nmCC+nfmanGWjIkOpHUKEhfRbqhkIh1ZXJGkzdoKr2Pf7oS
7oYKgo1C+FS5CIZThhxfGhVvB1rHiXfFS17WE4Pw+89d7/2Gb0Cf+iaKajjTHbIu
6YvQOHT4eO18ISnX8jLbH1dUiTkZw0x7IHM6/yq2RAaEpXID0k/+k4ofkM34CPCu
3H01gzfZmAI4LijVhKpb/M2bmaTushkN4bqyDDkLWpdZ7WEOfI3ysb8gWKtA/m9K
CG99zMQ3jLolT907TwWPGbppoh3Nyxn1gFQClLPgvN3b5Bbtp5kLiRC86KkmiExD
WdmMQxbP31jNm1rz/9g/Ziay8Gz4wp5DZ+2lJmF1Q9zF2ceLKl/Y2+u//1VZh5qN
h6bq52hGYtbdw3RvEyMNUPHykPBO8Nx/ZzsxGfKPlzgL53oT2MIcgPKfeLSbXlLc
KTCQLgj7+YvJQ6DED4zNJd2uC+GdIB87AiPdfBneWLH/trXFqde4gBWYAujOZQfR
yw/aB6hil01ulXZpl89GWFLHecI5BdQgwI8bZwl5YfZZIuxBqNnWoGGzh9UTudoG
8HXHoYgLJGUmCUUM3I0e0fphUstbTD/21U0cTGT3JECFk8MDdCRF4MstLXL4sHps
0JhROKlK8C6xxG2AsAT7HUNkIcU5vNsKz2EkMESMlfIgYnnGkwBVWDoTKSfnyXY4
W3AeoCXxNg8XnC35eGS28d54hsroSxHSnrLfjyDTmoEZMcUr8HtLyHJRE+FEPaDk
h34dhutrVYFOcMh5es67+wd5Zn1iL/4j3xMnfiR2zZGl/ljN0rx5tN5kvFNJIzXv
6+1xxHLGGrJSvgtBWye3r3hRWkD7zlkHeievsfKtlmpJhiP05Ug6dz3BYCmVOfah
MqaDmp7oX/E67FM+6RjU2qFdsHHmfNdZxn0rUdDeE7wrZRc35phLXPCk9IGdGFjY
71hnUVtpi/kh//C6F1I0kbXSAm4m6Y06hqtBUqOkZpvCmzzwGeLpTGt1iLDxqG6B
FLVNxAf5b/gt9ImV/qC9tGCYDCW0Wi4WTO/EVYLl0vanHaHwqgnNKhBHOwVpDgua
zqGhblxr9ntPqvPOOGPR1vCZe0DhjguK0xcBWCoYOmpyii3uKkDTpAw3St/Kz4Up
Suxut+/otttHWIOgEedA+lyOuRABRKVShDWnh0JJCgU509N0xwzuguPVk0l7hLH9
eBlMuGUABchdepvwlZiFVW6i0iqg/4phSkRKrqmtcIvnkubkOokMywgv2il/wc2V
+WU4LcExfq28dEQulRa31wwt9EMJgU6D86SrSEy3FyjgbEdsJryybe0mcOmY1yGW
R6Bye/J+Ms/fNGB3/hMhlsBMC32G9lKg02P7/jHJKGZXLLrRXgKaTq3XCFMgyBxT
O/Sxx40YZFVMDG8BNfEr2/kbIhtoilR4fWrBrcsR6iwypGWFWCXYjmrUMRfnFv01
tID486RXZWyoOVfOTn5jwffL4Dvz4V2uKcky1hk1CVxk7ueMeAzOyCEWKM9fXNbo
QE+5kmAIC4smyT39uam1/dzHQxGmXynlnhxVr7fpdQmeL61z3u8DhIvtN7mT865J
vb7Lin5/L5xln1GTVSkWIj+42jzf11njKYGfTadCu6EMa/Z75gLJsPliMBDwLVWH
WqxBbTAloFHinr+4SqoAmJlaec+/DTbQMd1i0qPJ+hSF95Wl30mSctqTohpS8jNa
wKAhnv81khP4vEMiuKnKhGo8w0+dY0bgSoP/osRkEgBi75KvJPxUrmxrbMdosvbR
csjyE1tGZgUo9XZbm2d3faLCShuSAf/zJ4y6Qt4vHsFGyex9kvSMN8zXh1PFrNAp
zswEmdl5hk0m4oBxcJ9lPrbr6GchDz66KVTjnH8D3QHGEVRW+Haw27QIG1U9lgMh
H4T7IQW7t+U7JUhk5pmWDkOv5wvJc9iRXSvQsoV3+Bd4EgjLVy9JfLNCDmhlmgu8
IIypJmXJTwItTK6O51z6d9SE/mu21Opcv8zvK3fu/VueyQ7K7zOZ+Ztp0bt8x4A0
4qHhv8WftmRxwaE4p9NgM0+d+PsYghy+7XhEgPXsdm928r4/PAxu/cgs1QN41+34
jeKZJx4dO2r+N8SyDxeejpGUgoXliL5/c9kUuw9zqpLP17ZXOjhZtC8VVcpAdVM1
4rSnlssSK/KapAJZa7pveSLXoT9u5m8u9SddR36CK9Y4zXDtaQsQFHiTxqhwUhpV
UxxL87I++/yTvNDY8ekrZv0m4M9oQJsUAwQAYdmh05epkyVD7b1WiIcvUAAnumwk
kduutLfNHAKtqp+VUTRwGL/5/atmWvh5yH8xEa0gDPUkOZkkRckf4uOhzovguLnO
lg+4OiJxEh0q+lQIN+eVTvOD9+yBrQwALM7YX2D31uxv1cXBMygkZGmnw3J5lYC6
zapWhxFEPYaD31x6m+DEEKb4rGM36yWhy6oO1sUUWl+tFvPP+//C8jZdPT/wHUxn
HaQ8Acr4lBva1JYCmN/Xj7iIJdRuCeIOs271xfdyQqid/bvGhroYgpA9GbRmMRUQ
3eICCyQDXzY4naS7oPgsz+fGsfyVea8mKORW3C9cs32safemtaoIk1mxNOh3a9wp
1s4agK9wmEyMSlzsVK4IWmqFg7Y6QmXOiDQaI5NxanfVjWPcPZj9pIqfXuHVZKDW
oCh4wNnBGHauiSzDl3M763gufzBo56gLRfKfMoJK0EjXqYXCS+MOW53/095n+GPf
/xjxqO12W9bPiGbXI5pk3nmLih9SlJQk2BiWBWTI2MhaPRodLSFNQaNCeqjtWr8r
2xQTqxGK6mAdaR1MszzKzKB2jz+hd7MQ1eg/2jVADgrex8tDZh0rRVF87+XVEVFf
NoXW+8iM8Oj5HN5oro0vUXzMi/86+xHirsOc8pVRsd5uB3Qq5la/tWKuFkvyarUA
bF2kVcIBB++flcVmVLg4S7a1zVVs1q0xcbekW1V9kG7HnPUTU2uMVrh/K7cPRut0
njpo/1jHQNBRs2wxxF7IwUJuChc5pWEImX+AYsyAu5303MW3DJpEIlfUyHNSzzZH
LE2tQmDf8964cSyxoNfI+DI8FDTn45h52SEBly+Z1QwaxCUTguboCIW0T7M3uGO5
rtyWcqeh92loYtxJbluRWSlg2WZA1EH2lwSTIWuD5Q4i1g5OcmsZuhSs3ORllX+i
Hz4lEd54wJgwCv9Q+EzO/j03bhheBtYgycGK+voAkkJqnwxxRm/R5i0WcX3vQedo
g5JkQ1WZQDIvhXgdZSMSTpTt3BUzzChzfRCRGE6NmOeY2KbSMk/A7r2RwymbgN9p
nVqHLkIEOCvlSB2yZZ2jJ5hsauebK+PEel2Am+6hei8+jxwCORtGinqoDyDMzeYG
l/e/qGxJJ1WBYQA48WZHDQsjQGQsX2QfZbWS03R44jJlRFQ/kqm2TWZvp0sWDSg2
GY00ixXGhz0/JJWcdNewZEVvevBZDn2PbiaNpzj9JSeAkLPwrK3rp3ExeCUSt7FQ
dyppQ2+HJFHJ9y7e7MHvQ3yDtH2B/nCEqRiAdXTq9J1NNqQU78sG1aSXoulzo1LB
joFf3cbvONHZQ44C5uvx00+8jM5AfBfF4So93avxqfLXCsatQ09FQ6Slwnej4yd9
fopsh5GfO3guWVNJWkIRArQtqNYjENkDD3QMhrUFOrwhh90OLv4cOmzpQq0nnwVd
HxQXOaw0dfdGwvmrOB/Bp3qxRkLGBJSWWRBDfdkBykVJ18imddmdd8ULWtocBW0I
kVPtU0csZt+nbquJCPWA5sgOa6WPjecOZc8Xr++rNgpYEYlGWBFCtntKCE+Bpvqc
nL49KC/GC3VACiONLbq7FezqjbRBQ3tloQMBeFdXfpzDS+sik3gQF1wEuWs5ZhjY
CFxwqbQy7gpSi5XCox4Nq5lbbODqmISOb/Xe5PTWjWVaGebyit43UYrgW0cGMNfa
LSquCOdoG51IVaFNA+eBc05Kav0gBeYE9DhgQgnzgheFM5Ua04UGlh4n9F1wP9Jr
D5rn+W8MGrCddky2uP+TDaPs0pcR3XmI+7crUmC992LMWUMEVOl8iv09C1uw0lXF
AzIeqH5T4UtzsPDWPg03FTQniWE9UQYfRSglI6LHrV/2y7zV0bwtMe6aE1EtLDpL
XZiiLnR9fVHYCsL8NDrjtxlB1YCxssHZyBQggcVy8pEYE8YXWZPuVLwZNTh3Q65g
bSlqBcbZ9Hd6AOnTvmZBH2qgvJiBmS+YsKquRW7OKn8dAZxanJoraVzHvitHcNMf
iKpH3OUFIvgiG//UfvB67AKN8Q2Y4XDo3xQtjpp0cNZSDXWfg3EzlwjZF/5LUWG3
SMpKa9xToyXr+iiCaGOSJo/WSeTDstRWjbIlINhIF8jgEIhS500kUwESdU9ceCja
agfi76MTgoljAksmoBCVuq+2+MCYcN64Dt9lFxMOiHfQFc4/ZLq9KwTvQBP/7Xdu
dXg6ngt1erd9WgB++Kk7pTKeLOaTyx9e/SkwrQSb1q23Jb0L9h9ny7bF0ZS2TCUL
8zFiGmVn+xIdsC/VOSO5snLsdwQZOe8qyfgw6Zw16RXyG/Vu4w+vQ1yaK1OEP4Wn
K9ooV3/zdgDxWFSDME6vHIP79WU2dLJhreBINBSO26IQYnYdFnpL7qhxuFena7//
Yge2i2OWArastDO48EUe/LSlxFlLLtwhoIN4uYKXzEZQGsSNrGjfihJJ2qXITodt
kgRUrPQ7P0tHRZwE1D92Uih+1w/UoKhT36RqaisxHMTVPrVOSAZuDTwWculSIZ0p
L2zAvD//ub/Mwuc59K2YzZv/pJBEg1DSa/Hz5EXOJ8617P/27K/ToqWE0/iX/84s
ZHLIf4newoL/X/4qia3YuLl39bJDJh6dAtrRADZt0FLhuRWIUJY49+AOXiD4ytGo
nBw4DEmOw3A8qcTVDQVBwzNYcesVHv4R7fOsSv4/hEvIVuzvJ7cWYFtWpfHqBuPX
r0t/yVwkL17fkFRnk1W/WRv1Mq723M5lNcYRvwhUQKuB5A9IiD6KO6HfE8Ezve9o
EQ4itesOWxGow5v7ufP17cgACtivxaID/+UvnBWRJxFGTZk/igUVOkRHEF7afDf3
1h4/0Kjid4YeLcmzLgInvSsUD5Ep78qy2Hr8v81qFfCotxuRf6P2mboHaIBgiD2r
ZWQt9jJd5DxP4jiiqTtx+TKkuhO7dNjWytp1ntKN69JiFlgxjkmi23INaN6cw2+z
fFuM3ulDFfd2vgVA+cnHX0wV7OALs9SN9UoQPHdjQgJtpyTXPE/33gn/pec7WQGj
HicCnju4NihRKm+1I8Zy8pgDtVQ5U9Dk1zdtoWhtXHgk2DKkULDkfbGQvl5uMWSK
sywmz1/cGhLW/P34rf3Aj2tYeM1uA2i9+0rdpWIEKLHetvbUEsvnNbRDRYvTpaxX
zMXar1RFNr2Ua/sMZspG/GgKp5ELQPZdWIA8hu9yvhPVODfaXu91fXsNShS4Awd3
d3XtU6ILOyyGfvHyzrdz45hLgqPdfMP5YGHcZ0AqI0EW4h3ocLa/70jWMeunwdQi
+P+cyIaNyvN1+qoHXeZMstRNXnHz8MJD4IYG/zTd25Q8urxVQwEMIaGRKbM5P1pp
ednOImQ+T+SjS/VPl/3x2czThI6Rt/h9tIYrKySHgthTIFiS7DSepTaLYKZZ7VBK
0MkIq+swyQV7Pu8k150rNBQVONoCE1Rx1fqMBZgiA91UHBeG43mDonel6lSMllQD
F8o0aefPSpdyteWvEc3Bb7l94ZTRBbNbOatkH+4Fw3ehU7lIO77im8Qzru1kswiD
k4DuQqJR+ZGwjbKnb1ZQ4HXxwAN4COr2e8goOKENux2kRS2biU/jXEmWc3c+Rqz0
/HVgulcPi3YrJzOu2hr0WpxTcOZrPuL9BZE7kxH+OR1f7G/jRJGSH4NJ6u4SRzTm
dTX/YoWYAFp5emxV6tkFZuOIgYr9IRhEcTjKmurrootrUYZK/sTZ4usPfVhmk2rz
LA+PKHvUq1Fiv7CWo4s2HJbC9I5Gc+WhJl6/Kp70pBsQOF4PI111lQ9o1EN3ZG5d
Xko4tTFmmXF8YP72SKcXYnHSIjgioR152A2Q9UqAMcKA5UCTKfTHLmeqnRhBSGUJ
ivatekvd8GR/GyUM+POU5ATydixrs84fS+hFKl+UtyC+tnmVGmUL5OSd+tjOeg5t
fOsVlXSmcvh4cyLroqeBbDQVE5VaHbrdU/97gYwLEsTFRwp5md0ARVvnBmdPBAbF
acjHSHzhBFDYDvC0hk8rwFuotr741rroQqFV98EcxU39QHwJE5L31uPn4qqgTTGz
XhYjym2oJAOyW7abxQvwOq1oRoKQCZmu/rPSTSXDIqnWKnG4Co3W9nREE4089ER+
45UEVLKg+REmhdcw3uJ7rtw4Id6ef2EpH2bgJn42+JAW95PwemUeVvaeI+JxSrn+
cb87lDjNWbV1DUtDwGCw4Bzj7QStTTpnsL5YrZ1xB5zvRfd0Sr3aTPliF8ZX+hMt
0hd1LEWJqiCQaFUxkWHP1+zn0OiQjKisioJ8T7WmFYnNFhqQJZRslexgWLx+1bgs
SxiFP6MMv/92nVMpQXiV0FGkK9Caw7Qj00Wz1zUx9z91Y/TnZj/PwSC0iDvMOyZv
bb7FbNCgtoMhfN9qMb9Co0XFYD35iYIHcpJJMTOai4hLdvCUjE3ZNil254fzg5DB
gOdiwzCZt+b5/Y/Yrgtye5DwVNn+2shi/5BJeSi0cATkmVljwTgM8OFLCXFdfBac
0AuQlMYzpxsIGRhlAj/cHCX1FAeNKSN9lnoRMTbu3JylcnoHzNG7DSswhMLUpB9D
KFd4p31lUQroWA9qgDqqaUZktKzWaBaNZPa8+8XHgvL04UwU3gDn2+DLMy/Dm0p6
mPNdbbAliOlg8TsFakndzb6i+D2hib/laQR1QHPmim3hN3+z99r8wV1zx99UuJN7
g759VzZJlezcvLmZjsXWasewJLsVnUp02vQOkUr0UKC5FqTUhEc7qV9RLayfrEm4
4gLJA5Fupzrh7PUfMsmCkxcF25/ORnxr7kmx5IBObpVFPZrUZfjc0qOziGI2m83d
m6316wPOW1B+o/MEv7kge8Ux7t3qukWUdnqpiDqzlBJo2i3h16c73XnKg0v7V+80
SBhCcigdy9KVkHbcSD+LBUCCH5+Li8cwu8tX8vyOVVj+i5dSUpG5PfxSIWe02k62
aISH6B80NZUdL6u5lWwCwUMQiLq5LPlNoWV27l7VHnJqUmsXdvzeMnxmUPhqO+W4
fF27nYfiYo6/iJG7zum7bsd9GBXaO2zEeeyKsYa0T/b2ErEshKHQ+i0hRV+nn2Hf
A0TuanLoyZfSpsWkzp22EpRQNR9BDTOJ7J5IFkgyQNZ7yA7qYAeX74Oge47vyZV9
vfRRR9nG5v4P1l1WT43cgUJsvtiEKtM0ko6gxI+O9Fv0PKwrjc2ARFXqWqeFwTtz
tsZhyOgItmykU9Vh19BrzTG3KhF9AtUihu64xjxxTA74k/3ANlB1Pfkm2XsbEZfp
0pKzMWIFZ6QLHQd6jTXXwYxZFNG5sBs9wC76LjQNxHs2SlZ+e07Itngdx3scGauf
fesz5aITwd+da3xClI6xGZNLGwaB3NWbctss21hiXC3MIccIRARcnCL1asA9BgBJ
81NJ7JjBB8Zt9zRuNUyD00nPO3hIBTeNJdB2L5c8u/U4HujZ+CRmddZIUiALSmfZ
jNIGRDwUKpoSX0y8JSbjXN16tC6CA3F2YzTZ852V1jEaFVt0rOHrVHGdUvXY3I7p
3lvuOACyQEUsJxtldvFDBLHRFkuDeodFkVD3yak94LDCXrnRstcLgjJY3qR8UsFW
yktz7bRaedQOl7VkE9l8RNxwpyFFA7HiR1sKNnmFnz3ldGgSmlkExcbBwntOlF4C
AqCBj4anevW+Yn9R6nM1SCgVVMusdq29kboUkvtvEzC9gErl2Am+BtJk9SkfpErm
ngjYrmCnXeNvKWGg1XEPNbLbyfi6DpyH7AmlbpXQPUty2s7SHm4HDY4D7rYkNVXl
dk9vyfUiMhpIEoXIf+HtqIA3TActEnpa1ldPBcUbuDoaDHbPqBt8JcR1mnSOLYp0
gXjCmCeNktbmJXs9w7OIt25buCU7laBKmScP2uuQasJWKtpGeRAkUkOzbf2P8zE0
lAcSaPSsdAXdVd4u2SSR288Akus8kzyg8GrvJ7+XibL9ZiUQVlRot+Xn5UWK8Jke
3d0QGz6JtPyzI0Z0c4a+A79eOPobCxD3eZ54g2EOxTQMhjjR2CTG0f31jcIcwhvj
9qvePi7iwjFcQTaKqTqeq693O647u0CbJK1FJ9/aYfPzq27jpHXhWeyRk/wLD/dX
otxbVDPQo50vMn6MF6O3DsCh0zL42cplrMzYdHHrBVDnZcm2ziEM9aG8v2c3ZOQ3
hJoaWrQl9UDJKtattkeLMic3FmOvsfHr9Fm3ph8ZpW1oUV4pxly2WfLzan9kWipq
uLZKcQyu0dA5WJLSQhWHEkmLvi6bbdlichfVspPez8/qpaJBG7g/qdJ0pJIqIYqx
A3Hjc81V84KJHeEIpD7ZckDcTsK+WmYirx0hlCj+M/J2B+xTEcE4oFzekOj1Ffnr
qV5LZA//4ymaxDSlnliwMUANLTgHmChN4WQSUUi2q6enXZN0YqjmUjTl/DbAfrxK
OOiH/RUs3941YYeWHHy+0IqnaWcaMy5aR8r1LTsEA5ck7slOTPV2kO0hFXEqGDlk
BMkPY8hEhnwTC8z1vQsDmpbGNZyURP21/i+lJMC5R5zbdflfZFkdz+59o0wn3U/f
O20STz8jYe4LfCPU0hpck15NMb/+caB7mczzJd7xhva0W4Qdn+y9pUST/YqZrfjm
6+0NGNQcQlpypkAPFINOLh5VUoHxD5JnCnKsximKJal+QpEAs4GqLy7GGHE974UL
DcPTA0sF1eSE5dSkLx/AVFpa8/2GC7m3t+xoQAPXJm9qgQH4nJ6bzUn0ZgI+1eMl
Jpid3YSuSoKrF3YNseT+0PLx/sBBmF5a/5wgCoEy4XLfxab93vYgV4BPbl7KdMag
v+eDOS+HU1m/xtd6S0uH6QiwyXR5ESwNcP9rcPsybAVuIVBj/6AwFiopEHJfYrYv
mvQ4XQHQ++Nlpwke9j6fTkaKLdbebvG9n8u2OJydCu06EPS4DSH2z61eIJL4kMuk
deXTSh0HQ7w7aXYbXagR4QKbrBewdXADG/EaxdIYonOzHxDFOYSIPdbx/OxJ4zvx
gYiBnWw716m4xok6zQlcqQxtpGe4i9f4e2nXju7lLY7sxdzMbkjVGouVbmnDfXdV
BJKa+sXxClFkb338rOjpFaMYovp0WKtm7EoiUB+OUTkySMM2wQXjBO7TvnH+JD0Q
QY589omRnU6RCOJax17efo96Ot5cBYOC2qkY1NOY7z6Z/ncPFXwtj/VK30JwBvK7
fkrhUiqZ5ivjFSD7DwSkVhefMlixmBd4Bc+32tQ4z7pK/zbs/UfRqqxzGpGrYlqF
smOKATr44jNUiMT3nSd0hVguGZcojJRdIS2ec/MgHbmPbK8zMajn4vUXXsYZnxIl
OiMS1jPZdP0mV2AIKakIPmMCpwEh/ZRX81eTkp86rZLFvAM8oh78rkEUdCe1rSeC
uk5gOPtP0xEkXDIv9di+/5dGZRO5Z3Q+5AfAoWC5qrNHLGOncd6ZxmRIu1Mn3v+M
C14LvDn7vbVrgEJs6nps4x9zA3mSgDvPrdW8DpZwdnIE7h1ffoIkThxy8w6XcCUZ
rIMZA/ovyZnzrIXnjOyjDcemfQVOXbOAZnQ3ZER9msdGFDXTe2VH7MVlkXzTgfHe
j8K+2r8ILBvjNSvFOBoE8O6TXGARNn7zdSZBjA1BnhEC8oFIRHWj1zy6wYyP2PVH
kYFuGTxl+yiYacPgpNZEeG0eegljti5UjNzpmFDMBxSyOaHuD/fvWc8dPHvy6PBu
XGqi4EgZLYWVyt5yn2XTbGty4bCm2ns40hOeHyf/p0gyZKN4KpjcYs16k+8g+EWc
qCfWRGXZdS1w0gSo+yC9wp3cHzX2HuoxKKiv9CkBckY4ZpSYgYmjGlRE6MxmX016
wMefFCjKrwqR9oflZNohN0DjXngiceUTHTXkxskmyRvJBCI0y6BMDHhI2I2CBl4G
YLFWvDJPXKvf3Ln62R/Sai2RHHUCfVerWUO6ZAg3suaqT8Cwu6HnqJRCe0Ozkjpi
YLCqQqhRwFfzqU/JX0aSn7MHLyG4797oOnHMvaANqjUjOhFi5pCq8hTG/jsLvLup
e6jkMFbcmm3zxvNLKWmiwk9y58oVgkMbKrImFWK65M2Jroxe1B8ND82FDYesnZ9q
p75/J+R9fgErtdiKIH83XRfAVew1gN9j2ne3hYO1btTE09WqlBrsKUc1Ei4hjaOE
byv9N9pnxXVXGlrUb8nfPHas4FIhhDVUekYNTs31lQRR31FA2m9Sy2DxicbY6WAj
tOcD6LsKncws63MftIfvTqwZt+8joGqtCKxKW7cIgQlz6w9CKshXhQ7tTpctTPlh
xMJLYqZyXc2CkhIMraKBD2Jw0j2ZueBt2BnfyFc4IX8S96aZErjDCbBMrJ4P0v2C
lpHJ/YinlWDgeunaoKT5kWzHMNKGz2Ihqj6F5X1s+zistq+BRG2eUv5lJ4D1svhh
GCUB2Mswsdb0jGDEgmihtfJI0j9unaFLDmTLz9+6awlZiL/3a5m8dl78+Yu+xQFi
PXlZNNl0xDCBdSyQZp/NqXVYNTWVvklC/5gab9wYLpEp1FWY+KVQjO1I//c0Dl+J
Cwi8Q9M4Ml4QMSzbKKGCBfRkZAcHlGb6y5bZDhOAmmeZL5up+o3jPltt5M+ZQB/j
k19tfzA1oZh6x+qytKoeQAx2bGDCq7stcPHJ75MPM9SastJg6XroV5mVmRiS9DIt
aq7suCr7i/HidNN2ZrjRoqqjSqmKbc4v4L8ZfuSnL54eLv+569TTsPNCwHUos7wD
z8wNVWTnFR3EQ2OEeKDopsyY2AyBQcamZLWOvY1DjQrGqFJBKBuW2I6eciiKNbUg
JK/5SmU4aqYXsevcY4TCJsklz1cHNfI+iGk1bbct/+RIw/fZHm2Y098knalMAPmY
61Vx/RPEsL51HSQDGcXKQl1egpa3IHB5Pbhj/xXsJ18ircotLFNCWoNM7cL95yIU
i1lvBKyXsccRPi25wDZsXvzRraCBH+98SQ6yPoKe9PlbbobTHrF2IheFNDhnsTuV
LNbBj8FVzpYPhfJxtZYHyNC1Wgm/8jmR1HvPJhLEGbMRHBb4wBpYNHNCjlLU/dTV
72ic+hZriLtDSBTx5tmhJl93S6n2d74q6sQK3yXiQvHI5Cf5pqbDcSsrHewV10lh
dnpAsHzOK7Yrjjs/82VbGwHqKslwdNHpzbX12zmbVSkxvBWoy8LEuOyT/ntpCvLY
Xirk0rw6mik5N2LKl6HWyD9OAPDr/r3kjN13FRuG+IicesX3mIBl2T96VdjSPcve
iqn8TAH1dwAzVe5mlEXdHxxDtap2PELRMAncwbcuYKU5MiDp3LGwqChkrWJ6AFxO
B1P+JhtJRF4ka31+r9nDiXsY73mNfhhCwylPM+k9YZnxhyvaiMI2mAXeBLJUmx1T
Gf9z4bCaSxsXakO/72D1yCv3SmUH3eFYusuPqn9Tlb9hKYbXcK7YSeKqgQ5CLPiP
fylz9KrhAyQxPjaQbMAP75+ulcmkBVysMwKactdL7QPVbwOMSHl9wEL2DM9Ktycc
FEbhPlVtfU6SjUwIzTDvGD7kpJNa3sAmzy58qeJujTIamUD8V/UVRVlxpQ3MB5f2
97YqVr5/Geq91iWVX1mDn9GOjmE+xUN9y4RJywjmlm2XDsMlJ5l2zfWtMo5I2p5p
nH+E5+6yssx/ui1ZMm7n4PQxQMrXVAVQfMJj1CpLz6UEU8s2wkBY7g+SWKrCiflY
uIcXIvYL/Lt5EFsXAK6rTdS8IWCmb1sAcVPs71BeEVIH4u/SSlsPbKKPWOo9xu7G
wvUlrmem5xtv4MLCF6tNiBaw36EWQ9kkb7VsKNNJi8Iy71fXAYNRtBt/Vv5ULfFc
qpw2UUX8Dxur1Np/YA81akegGAk8BPvq7Q9EzUOzaiNlnkFuJg72YXPjS4ABAX8y
P40z/luCvq/sf8RDsQOVwBs/+HacPrpIoR9UD92kMLjyF/hSPPpBYfMl47XZgutm
feP8SCzWpbf3yPsAlmqDg1BR9easDQFVwFJfUret6j4a6x8NXsILDwi+7+TBEdID
41aZYT+gV9IM/kdRW+mrghBVP47jFKduKeGuA5uKdj4GBhn2j9FzRPKRL2PLgWIJ
dUjfpB0o7bc1PYP0KO5jcdc1nWuqINwOwlPd22B7HtVWRQsXwm23MjQ1Qgs0dfjz
znf925GFBrfvuoPL6dyKjrutsuVSW9eCxylWzlyBN5Ai/pa3niGochAlfBTOMwez
Z7OliqDquPlyKJDu6B0ENPNtKtA1as8PH61mUbtPTTtSmZPw5ispkCOYPxQpmchy
3mBZgS9WvKqG454WxOV9vMsl3eTA6e4nFabvZlT3vGC7wyc7uSzNZC8e+gHZotVV
we9fjlInTXvI2pA7TBq1c42M2aamIIPk0noS/iJZ/8YBzUdnCZPIbu3Q2QSPdlH/
idDiTWV2RAFFEoRzSHDmbVZm5GQ5ao7DeyvkWFXXZI2jsFx7jusieKNGaoFvp8mq
wjaWBFElXz4foZp2RRU0MRlGrzV+PNQdZWpqCXqcXMwsAOSDtje2ODo96ECF+rfI
wpMMDKspODWIMKBi9NZqXPRnFRc81tM8Q2pnaGpJAMGjpk8R/xUtYMcRlYqOg9DJ
Aa4mDB+kdnu2w1cx8VZAWZHFn5pzdw95By+zgUEEYEuBra+dF2+vOzUyZhGKxN7+
0GZ9odWmluFiuOonRexCnUC8pzfmpNmniltHpQLYThwRt9OL/KL4eIiyqm21D40f
8U9cpagZKuBxjtJqSBLE6QKHpRgpU3mn+VwDWmS3UTXzBvrE/qev9PBAqQpLo3HM
U24ZLf8hl4WaqAApcyd73PHG79wDY/57pN1h/jcnZtxD1r+mW7EzZNYIyiqCA6Zd
FAUPGOlfqsmMO1/fiaicp4c2RyMuVKpYnGe05PWAi9tUrWn/2UtIH9QNMhvGZtrr
pDWumFTMLsgIHuLq5On0E3/F36tBbjB54of4mpItjw6jqsxTOH185Vkts8Ot9uKO
9k0HG4lAijOgB5MiA8mS6ofkYciSdq1QMp0zWBT3TzuS3p/34CZulRPN1zA+Hrsv
1kkN082R7N0FE5fBvIE3qQEIQcMAlWfs30AiTaVL2GMBUOOFSy0y+xgSnXD7nQYl
uowv9S0Tprzb2vYn80scghYKoh0U+y6Qd2W+Glyf/fvrh4UvqYxPvbM9HL2AUEy6
Uk6BHvcTphAaYzjAdVXau9ktpUJINXrNOv+CkvfoOV1jeFAm9XUImN9x/Nfy4gwb
/m5fT6NurJNFMUsO3D1xEGxi/+r+YBkn6oSt201IUanJxMPp2SSWtHxAz/ua7alE
tqrj6SymhHoJsLZQ/HMui0fGau8E4feG2nJMHzoeTxx7/Mi0xsBwjLqMKuhB5lEi
Hwt3rP34pQ6s3JuWG6Qbmxq1KOxpo+Wp8pItA993EVOGNLj29RsVOgmBsd+shykI
Q63+ODnKTuhGjM/d4//BEqhhvQEbbhrus8NLqTMW7DFWVBGGpKctfMi47ksWOlzV
MFpVmAJ4I6Iv8lxNtlq8PLtaRaTAMDkpMS2nQ9QxpWT/fyEx+Eu5RbEmo/4+fRSm
Pj4CvgGI1UI2VlQUkbqv8jHeqb6lTMyg5P4NXJqJjRn9x5IsEhIk8gO9ttysUPQo
g4XZNALG8lv/ano4WxN7/6jUFTgZpA0tMaJb4AAL/T/pq1gMjA7pJTh1SlA6azfF
MHLabANqzMPe+Pdyrmo8UIS24vsmiajB+DFBKmS0xG5zzdLYZ1d1aytKb9/UgzfU
YrJmRRCfJoTKXL/q1lYvIt48qzzi4Nqm57kZFOurxqJFP80D4PQI1T8rncikBepy
kU+JwHe6h8udW/MpVFVEWJnslht1meVIu0E1KV62hAhasR30LQQxAJ4vOvuRfinF
9ZyIblnAilJAzwXoAZLVEAgtxGc1RkY+G4GN5y/ugntZH9CypMF30aj0hzoiRYM6
vgHn/ORbb0ZhofgVJs/O7NrqD12BNzZE9y31dcOrVO30lunaC50YK9yAvRGevKsO
4NQX3fihrYLkSiY81OTAz7Z489B7i/OqsBKl0vc9M54NY8624emWRwZfI3xktO8o
kzYhensk6c4Hvmb86hcZ/C/5PMk3QYfftxEymrKUrVyc6J6mUX6W2NBZyCnirejC
inSrPR3yHwDzZdHXXjgALgZWJPn6kTh4eErM46n+V2mV7NWgsgzGBYzbxCAxfqyc
J2L7UZSy58Hm2qCEn7M671Qjwwo09rh9kb6eV+HOErvO/sqV85KChx6qNOV0W6zA
bgVXpF7EaydqCqF+2y0b9IsIkEMnfWaAwd0KtASjLXmojroq2h0d3eRROZVXfrMp
8PJarJTJkHSxcmd1d5uFXoznPNJQSCkBNT9gxbkr1fWm27U8SThRbWwoE1gnTURI
zgBh+lLfy2N+dU+vr3f6Ys5YLiWcffZ78YmLUT5nk8f8cNohAEjrDRLQh4qmlpbS
+HPGXi/uHLQz6OMTyh+H5BTIW+ZU93AGKbwqmeLsvfLSRzTjij6dFtuQF6ASQ2J0
qkyovSgtZY0EdpsrV2dld9PfPFy2W+XMqxbaBT5kYNGdUhE60fF3DJiY9mTfjFrs
YDXkmUHEh4pc+OjXkizKjmWVAWKs4um9OicIDmG8ijqZOxoanl9KB7ktYvz8fXLh
AaX/CymUZZqUZvO9SQ116jhOU6F73WulBa8B3BGIsW+WFXHTku86Ot4Xr4gU85Eq
Wgj8+GnYfTK5grqmP3mNCvXKDg/3zYJZPp0w1rCWa+ARmnhGWog4z92ytofPa8lQ
9dxdvfomT37CVz7uHvdkyg6x4ooIEETZQCreJdBnhXPbZhBG0fiLNl1arj0tXSC4
55tzASDMA5TN823n46zFDiaVAnXVcpbIn5uF0D6lmbcUZ6SHKCILBkOu4bwi8Ok8
ra+oApT0b0896au1im9AqeVI2YrP6iz/0qQwXNBr1LT+WFy9YrGDnV6TkyG08nzH
N9bxpJ4voblZdvh81MXb3rS7pZVuG7AnHp8zWoyyHTszdK6Sf4KaY8EgB+yewp/v
6Iu4dWEN8GOh9wqLCnJNY3d53GzQN7K0ju+x11U6tgH3iZA8lb4kdEY9R3D/IGxX
zDwO2slcHlEUXAZl7OHNoB7RTqqAsS+0r3yFYsjYOpGBVmeGEBdbdqnuIoe91Cd2
fuKeggs04MibCaJ3nlOMX8f1kM+ZWf8FwUn1TSwI7ulvjcg0doLh64SsHyLO+vo0
+8iK9uSz162y7EKt0IXFayS6GDXgYUFcxPCcbX1rCkbhoSDGJyoWP7+AfHYa5MMf
DbhnnZv5cvO3dwW/mOxZZRSUKsuaPVPZzZHd898uIhjuenb9TAYbSPm/GxREFc+f
SnB7upBO5VVu9W1unQuHclFiCLmuJAm1k/Jo/kOLTYh75nW5khbaxCB7F5vgG4ox
CDQ2TgZUDQets2dOxNrZ1GOsc62MZXR67DuW5wxvY+UrztHK9LamB9baU75RoXL9
1aBmQ+m0J3raCutpnLkdVZ8vzF1SvYr7sRhfdGWkBgIUwleJhQRP+DhTl1xW2zhB
FlhRUsuiHw2usbjKav0w+Yh12M4qYT4SCbnzm6ZWQo6sUMmvTiNUDE/GrNfrspsk
JkDyQGtTbaLeSQWyKQZE82uaSuvxPoTH4r0fWFwbSofV4NMDQm8iE58UKcs2crtu
Dn6GT0v17soFcmrVY/p1ZdLZjaAgkWdxgeytW150CNGaechKkn4yOeIUFRgmdr41
R+z8ei0E/RVOkSeg38Qk0vjoO3vz0TVV3z+XvW3x9zsM7edGTU4lmcQXp5UbAIZt
yEfY71JTBDh2N0NfHxUDUzju/upOQ3J+yhOBvf/kWjOINTmc1EuHEtx6Ktz0jc22
77ExviJnWugRGniUJMlUdyXdvTAjGOy5QRDzEWWGD9XhQtgmuH42yJ+Y2RFjQwFY
mp+6tgD8h+6rLa5H3U4o212YHv8e7xpMS5FOpWwqZx1KHYYRA8D5ZUHm/07DyQsY
V3Q5nkXhmMIgJ108354SUsiKc+tNlSc+wm8TohoB1lXEdNFlOLxMZk2r6tgptLLo
d8N78rYf+lY0LV4uifaLapANSZjddwQlfjc31Av1xeF2s1dUE1UGLvDEfWDfqvX4
YF06MTG55XltvMD1Ik8xdpti9t8Sx/tEuY8LHZJss9kdOv9Qx+g4Op901Gv5JGWv
hT0w+1dqyLw1ovy2djC+EdzvLmIvUqveq1C8Fs6nsdHId0icZDc9T0g6NVxo8EVm
oXvhkL6BZ//hTnGbHssMolIGFx+yGA9aZFkMbyzxZ0MSPRfiL0x8bMpMdKpl6TKh
fasLIwhA0vKBKUr8Z2XFaGPTSfua2CmQyn9SiuXFIft0VUA7QNsb1tij7ouwknvz
L4feRLlgbTbvTyDuR3KaB82UJdielI19K8rDErJm/GhJNZj5LguSF/lLVJUQMEn+
6LzyKIPZsvDNd05dFQChfz7OueuVFQVSTnplLHoSn+pTr3q0y04GYDCH3hZClY4e
BdaEj7+X8uEhRicNziIECa7MgsfcsXbirLL2AJ3sKUKONEcvsW4r9ffQNehtqee3
GFI0qiJTtLbWMxihtTpldolk1gtTfc7vMpEUQy8VCCNlDF5zb0f1Zm/KVnDxWx2T
YfTo8KWEun4+w9fBLvFZEedqR33RJc+BhEDl3bSNiCrmtalyIpwnzyK/hOuKuczt
43063dAy8cfSi9FpQEkxv4gL0ZERTbhA+U7wwyY/HN/AOytz5+CA3XTrXh6YjpmD
XnLkY+BWQpFla6gXy9o5sRG5HusSR7HQyNW6QKpRZq9al+n+kcKjdciTvAhF2zL5
qrmJxq6SdXSdoSXGCMGIR/9K0wQ93Fig6asPENqXzNDxRmbUDUcSgSY6GJalSCOp
gbcSMR8Jwy0c5tE6AqPUC9M7lBP2HAPgL2QrKaka3qj5PJrJw6+VIgr1APJdkxAM
1NxiGrtgiRiiYeTG737TLU/r8FRW3nHJyJWneAa1xM6bC93GszdrUwrEV5iGBSEl
OGYq3v5RnDO1LWWEYMlgXX+jKEoiUlwzJ9W1xCKkPJIOOuC31bHZXANl80goJJh9
Q2Owse9CZ/iwYlz3UJhPMV31P7FhQnGhOdPb35NVRq1QZXMKTc7ziz5OIAEarmb5
kCim9C4q9ihI/2GaQWIuN6azZ5EjkOlwkYK1UtDNv2s8SSKFPPy5F/pUzVdt/7pI
bAMczlcA55CkdgWe+L2Mlf73R/wj3IYr/FVUfF2m15mPOaOfSXPS0RcFxWLWk1HC
Buw+ZaI/COfK95xeZRLEOzu1f/VqKqoe0b8p5g8uLB6ibgKZdalGSJOEycfdkwcs
Z66CmR2dw8PKHaTlXuvc0YNQ8p0JsUdTKUQnnAifKwfixLtmIoofDVsfoZAkxPaV
Xoe5XJv8cdwc+7M0gyIt6V1guLyWEiFn3MgcdafbrW1q5hEK6rclg47MgUdhNc5v
tv62FV20Ln1PN0Ut17D/hw4hAMlwhurReyNVmuKn06xewlJqfNxsmEV1fu86jUZM
gQyEgjn668YjBAaBnn2HUcS8NRvmRTY0P/khDWT6jo+q2K1UqomHp/71au9tBoiO
/MerO7kTljGnpRdcbPSfUZlSDcRCOEJ/FBPHsGKFKKpNdX6edDabHbHSHCuYKG5m
l3qQfMOTyAZo7A3XHJBPUHOOJ2bEODo18dKtw1eQTXwPjgwnzGnt1RhxLGwXMmXa
bqEVXK1utb+a1t26fojwvt6aUs3yJba6+OQB3/OvcQdBgFnWrv92CzlO8RdmuWWH
K+B+D2o33oTnTeY/YnCH2+hgW3epsjq9FUwSsXr2/j3p2pDr5zwxbH6kPwEzVRSM
EEvk54CY7pdmNZ5sfE6a0FCoJlC75nu+3nb6kuUex3UdXpRw6pt4BQJBW7XaVBrN
aUqLLtvrZvI0vrNMpSGqwCb+3trui7S3W22nzFVCfk3OmP1iSClgLz7m5XQwi6AM
T1jyFrKl1hO0AmWqSPSH7uMGc0U4rpjSGJk+rUO+F7X9qODIFN5ePFqJeXnhSAZ3
VEswhdWmBrNhhBUkiuHipF0FCOyNpI71HKLXvfgu4h4KKQgGpk5nohoyFtSKPmCx
k/4ZkaFIBikL2NYs0pTvG7PDahU6D/HBzAcwFLfM34sZzO/hJXd0Fz+ahK3ZmQXS
SorS1fVPgpgKas+XV+z/+iZbatsymlzhL9iHWt7mx9MGJKxfiyQ+RaOKDzqEEfCq
GTYcYvJaJa43S+U0tsSmgG43J/zKl3bjuUN4U7vjC0mgKc5fQ0OLUZvAZuRjfLsM
5myz0GsTIWibC1WBMda9ciAjt+uEwYPTvlPsCHaGo4NVdllX1ZhgMr0g5WwSccPm
x2/fvrMYO1zBnvMEK1NVhCggZEPisGeJuDoqy4gIyiloRDfcxfQy+D1LsuQCbCsH
wnrLPtDwc/3+OhDCCunDnUMuEsbWFV/4xF/HMDnH72/DD7j2c/ojSnL3WJlZXnuo
oTmLG29oSzMfvMQIqLsIFskXGY6Gt64+0lzKfpyj/k1wlMtaEgKyekCb6yBC+76f
s46Mu64VKlP55hG9Raiky4fqswCbSUGaixq7pF+cWiSeOf2+zBYgQwDZhOsaDRXb
N3X0LstKHljkhBRzRnhhD0J5Vt9n1Bw2F3njC9Q91NMbfvydeFCw0dq8TSZiV3ab
u2kBC9XNToJRplgUT56e1HAikF0nS5jr/kcmd5KIZcEAj3d3x7oGevY3VFOuI6Uk
4gUPCYYC55tWMreKO3sXLAp6+8v/JNmhXWJUacoOaUhEkuvoJAegAP+KlHTI+Cpi
vy4UIhOCRBh6wk7VmswkPdWArRGsBQv1Y6muX3nMq883yjA/c1ymUwDAjb5/Ywkq
pPdDRADb28fpy5Pl80VkvfkIjL5oJXo8Akp0YlDnI0tuLrbG71QO87CScwEyhCWv
ouIkVoyEhj+Xcd9YncmOgGTuA8aEdJCr9x9Ao3BBAfIczU0Znuz5F05GLBxmZn3c
9SeDe8K7/TNMh7avBGkkboZz8BCf6md2og9fUT6M1n/vXyAIyJeVV9Fbjwo6ap2Q
AO6ClDoOeORzMEIRQDe2ZAAauwvXhMQ4rAv7CZ/tIzfOGTmmFfRJimKOwLu0aljF
r+3K17jugyzeFHROQc0zkZuUs36IPhG76q1nztZAF3cbiAvMJUZvd/BmAgY7cd7r
Jtznhq3J44lcNYjkEl+AVQv/znePWA7GlGcvb3Nd35J1r7XuFV2mnKiWsLDtgU2m
RuRa5N3mv20c6SEEgYLLcaknrFeuIhFljCHbAYhK2PKiWtxRwI9FFy64Z54ScmCZ
3Qb7EEqmeo7wAA7j2mZkphir3QTuJUkUwEUfKgkDrKl5mdvd3Un00NbXNcrG+jVW
reMsDzrNtIfQKayRrAybTp6AViiNmSUKopSKdqBJEb3ar9LKs1Sxz81f2dzqDAYE
mN5sTJ27pJ2XCnYgCkQsNqHQiVxx1Rnix0r6DKtioUBA43GadQ4nY1DLDRQPDHm3
JbWYu3/a6dVE560kSXYwn1PTlJ0TyRFO6Y/92jKOCLnQsicz/2nZv41IBllvZ6xa
AN6ECmUOGBb4FrqReFtFtKmFnyQrTfrS76qBO15CWv5QWiRgXi2NnB+fgIvljF8P
VM7l1W5DsZCp9UY6qu5RHboH4M9E92H8i11/nh0STYSUBEKaYd/ZEvFcIVKA6Ypc
8Eobu8a5rytjs2/KUVptckq8mYn3H+mi5GhlfQX2kNZJxRJOLB8qWhxvuESwHzPv
OwzkMHiguWOU5KrJZPMCf1Vel8JeykGqnuqMFUoE5kMRYxD2CIQJFFRDJtaTHPZz
JNFYAZiS39nVSrGcoi6ukta3FYQy9zYvod7NltuqiBChJ80l72t8mtuVqFhFytAs
L2NpqWC//m97xzyX04mLXXkgwjLR76fmDXj5tXTHa3YfxWyh8Tqbn9VksJa+l8h5
iGv29F6uGtZ99Y9qhRSl0C+x45xOoffmbM4yHvDQ7GIgOcAn0lzN40d2JMasFKOz
ADcjYDvnvCgZXUT6YJkoZw7mnNks/6z5wqVc0MzX9XWyRAf6hJhMRz7BuHlS01Jv
AoznLHi8dmm75z0RNV2HSFO5CFpfZQUfgkjvAa6q1R6w4CCXPxBqDLnp5wvDwmi0
a6qxnd2nR3+VzspXmC2rAV/BLruzWthfs3BQHajRMluwUvpqDmlsQP28eXg0w5V+
KmJGNF/ROHmkbiUmdqoYXTtSQ84H522iVAkM96jkfZh3lew4vBfoAd6AOyiLmX0B
U2xwrw+FPKVDwp2TZaHwWQZip0Lf2KtC4lEBj1/XpxzjXgpAZQKUsxuxMX0N6sW0
ZOc1VL/h/XzWcN+0lb2VTBCQTlUTNc631UqrCkhI9/QIYdoRHM/335mPtgSKncf1
gCHiS09871DgtYJwp2xlEpCDapDKeN9Zt7F96SOCsyb9y/S1jumqeUxoUBzkWVyK
NaVPlrG1pGdgXRucuX1epx/ofdWUJDVFLjBM3VlKtLwgiEbA3LtZygGTSi1UxahC
K9+J1a5qyM2666780cLg2chvVoNvBfJ1fAj4hjlLAJ5sE3dg6IQxSta5wLA57Pci
ggjEwdpo6yvhMsoQ/AgtnBwP6BZWloxktqrd+aIeXjKLJSvFt/SxRe/BaQyQNc4S
7/bS9ZkR8BVszR7zvzLFDcup5u7s+QwEui1XF8iXyBwf3vxmsrQwwCqlTdOVeKxh
8brbzTwdjpAsCUqS190ADsQKm3xZAeaZw6qgU0bZcJJFiBMccuhhP3fJcnoY/knR
bLiL4JrUxnl/xaN1fFx6IR9hMynILk3dJ7P+wcVKk+QFPvKK0IocVkDQ8sN9Tyxl
tpMsc0tgWXscBONxThNg65pFD7n2aVZIWaR5hRyWX0SZs2fB7iV3c/Nm0+pYbyAi
taaBHFcN90g4pW3UpIC5b7dcgzw09UhjMEXZDNNRAGIaiYe4KQ4+V0hOFr30gdRA
4Ah0p9M06zKv8QSFinh2gd3bA147XXO4LC2Vpa9yBYmJLZg/BPLfm1wGrhi4jQ66
Mb4j98YvdWwqBriunNso/K5EMoNv9muaRdFstvN3OpWdpyD4tVjHLJ/BDIi4/Rpt
ofVsZqn9ULOox2Djab+SFA1T9b3B08NjNGLcZj62dGSWU7USB7JsJW+gJb7QNP9q
dqwu+7MaeUyqfs76n/13pcnQDWvnvM5IVYrd03Z4d4uy0DZ0vIrfXIxrHi1UlwK6
YJpOiwv3nNBDvIMgnsQZ6lujlF/I5PK2IIW/iUPdNcKD5wCbTPjR7jG7KE7sOVRK
k8w3D+ziiZC+qRlo/BJQtQprl8mJVJIleI2HJO5j0gq0po0DwggHPF+Vjpo3xFy8
V0K5A7o29/m6QXWamd9mnaQkVMlNmoD8mv7+Zhn/UKI+UsvZQj4E4k46AfRT+nvD
a6vdvg5Lt/ZL6I/kMiNA3Lv3TdKK23cvEUgWyp0FUgXV9szDrjVuJtjmE47MAGla
ppgNbddqQNtvzaPfg0zFvhm0O+AtwRwz6Rmq5hY6PDEx3yaMle+pqIf2LY3LRRdR
EYsAOVL1pNA2RIiJzB7Ii1r02yjc44HfAkxxdgNO9H47GVsfs340cj/bJhw+segm
D92u7PyVcbq635Qct3CHxR+lX2o6SsXtOoWmfKMNpwMQq6vrR/XtD5OEbnisWAi4
PIDcIQg+Mh+DyqLfdOYEUdstm7djumlaCPZq30tuPJh0OJEQ7RvvBDoi++wvARGf
HM3X5lDNbfuKHq5XLXVtzE1wQJ5S2kBuxMPJHAphb9SAc5g9YxwigIlT8rovcTJi
MDBjo5Hj3yN/MYJwXryRLwJt/eke5M/0XM4jXT6+Fp9zgBEOrkzqJcmK5V7O7LIB
EHFm9bSo9x8cGS43qNKyFeLqSqwaW4Gs44fzWIB+WQDTmZ2I69mK8F5gJZHDIQJf
URCuzzZBJp77+s1Hxh0L3rly5opkFEHnunTGDWKQX8Z1PcbsOOfGiTlNiOCg7q8A
7aZELWZBH8uc/qy+SBFuRMd6jvjn4Yk0jMphtVLCvwg/rbDkiTXE8KdILbgQX3vM
mT+1vLi4HboGBMRUDxkkU7ZO68jMvQqFjF/kYC8r0Kz0sIprOGlrJbhm3WzH+UB1
Y2TzpEGOHOpcYLzJTw5jsqSiIrQEdK44eYWdahRJvIfCIaWWAm91TlokRY7+UhnG
xIIFSX2uhvWp6Iju/YaBZMPtbqC5X6EYVBM/nOLdxuECiKzPz4U4bFBOxyAK6VSB
pQx0A14W5UI9m6EYFbkkmWP/up8ca89wnv53FRgGxjBAVqxK+fCylONxwxRlvnAl
Aopn0SoAK3u++flnDD2y28wIC+mM3bKfFNDBh0OC+bHnDdMcrxIbqm09RJ0/Qxo9
3CbLCwVmdMtzpTHgjP4DsUOWVez/DUvSTOSxBddCirYi0tNK23cOaa6mubmRQkU8
MRLZSqC6hUdmwBSze6U/Ja4GjzFNmifV2vlntlYlFCa4QfEJ6qL3yj4Bbx5k+Vn7
FtWS+FjKicqBAkRxw0tQK4EwgRAGnc6JUEPeaP9VS7rrLyHaoss0tQ2LzLSiS41+
kkE6jvuU7eVSiNDstnXv8PMG0tY5vaX/eO36D1oV2aoJmmqHSjrsTTJtVtzJ8rNX
I2ivHhxf+A0oMk8Vv/hAJe5zIydt6qt0OAoMzELfNviYZQmITsO+TWpUANWvLXpM
B1aQGaL8OCUMQgg0cgMZA3LemwOI3Ow9AYH+F/L7adDARAxjmSY4JuhoNKRzJznV
Zgms469Xi4dBHy2wk1ZJFhJk1aIZi2JRFS8SwSAX9rW7UK1B27OFmqWe73397CRf
ZXZCvxdW49tKCZYuMHgqn7eDXbePPPcTwkvQw8Uh7/0/Q+Fr+4r9ZDEK/AGAdHfZ
kqk3/NDL2E3NMGCm5vD0XaJAEAJyLqcUi2+TuV/7O2IEJrxDzrHJzlBpeM59Eaky
qIVx8IKchaAcmUU7WSuCpWGbl2FlIB+62PE8Pmfr/n73NDjWfl+sStWCWDOKRtoh
yhGUpu8AWd8Nf9wgGXY21kU/nNTvqYuoGTOHoruFUJEZcLW8BEAGZytXeFDE7494
t4Rz/Ia9sHZx8B1VNbwNuGjFVKu6ydFjqKsTx3/E0RQBH5lnl239rApArOAmOpBA
4XrbX249Iv56J6qJZS7OQ0n10M95uKYYP1PQhyrOfI0AfwnQTPWtiThLITUZPy1i
/n3xicCf5XUIQLrdDFRp05TbUoi35ei1ClUpHQxwBylr9mFMLnAmgZhtMFakGNjr
y3tOCMdZwdBoMra/2Gco8rVUgaqCgZdput7dNz72QDBLfLS8uW1fnDEzWNdOd4Vw
CNJekV53bZB08X/Vafoi061vGOGu+D+WtbkyEpRF5MHAyzSFvADNebUOSAZG1RAK
5UzbDDGbssbW/VuuTiNMNl0AUKUhWF3QZwDolvhVXFxzo6bUyRX8TaOMG17S21J/
GTSieWVyVvbnmoQfwuBcVfpFfLr/+HgT7KV/sywnfNvXcQnXCvLNFVAeVIecmymz
WGgzp9PcXDs3ogdcZhDIvlxKIwMe4ee0vNwj+uxDH0PB/MzUxJHZqgg82gB92FUE
qYtVXT7jSAC3toL79R/I9ig1ptyonnDrt1SA1AETt41AdTfDb+WkoIu6zUZkHujs
zb2txRxBDMDMl41QgVDitaBWXKfROWAC/jdonfpI5ViLYN3X1+sINHcf918zQ9Fa
EPO12xwC5hfTPAVlWi6GT7MdHyYmulJRiPGnm5d3zo/Np419nK/UjIDlHYsp0TH0
kvm+XirDu7lsLhwaxNL0v9ZvgWMn9eo6G5LS3nqkS0W7P6BDBjvifnNZR+sRSQUA
MdZlquUa47qt1Nr4VgasY+eek6Kh/IdIPyl5VN6WKkXO5ay82SlyAp2kecrU0Vk/
DhyI6t12KdthQM1U3fO49MRow7Iu8RioXqFcDlEdrGfPL9Vdyfw4xfwUlTrmbfOt
bL+gQbOTdhgdg66OUFSUwos++wv3zz75cYBkTc5SWF2Pk3aljwrwEfcwt3oA7iVI
DzVFszeoWsliGk+Aymta7s68z/9rJGSzspgcudwzQH8gcBM4LKRAm7pITGmy1XRf
7/Nu3izH3cZosisGqjjxu79l8+ORfK5sC2ZhasiltFbZ+dxeu99HAF5xGJXRFEqC
hA0uoeyZPMYFvHuWDZUWHubssLRtd9wIqHlp6008WRNsQz56CsUxF3WQX9Di2IPE
oVECAxL0cPoqx/z/iLYTrGTA4zQAg0k773n2U7OwbbYw4W6Kdi/ZHTn62Jhkc7Xs
1izqKjdtsDnKWpdWZvcnq5xE3UilBLgLmpXEfQDlflTB/FmestYVQBtUTIQeCSpJ
QUNyfbqtw6VSGmF+HfISFW6f3ChF3ZzonZmTmlbBwUBlRo7aAWE4/+TDjzwoUTcb
A4WYiacEzLxsXOTjWACdgG1GwuUF/5uFUiJQgPFFISUBhGptnKGJM5NXX4t4utK0
uHfg9Hx0eEe/Lqo5ZSnEoHTBM/sug56uggeZ3WwpYynBGzetHhqd+jRZrONOKaFZ
a61BL1rRv3d7+NHNpAsjKZFAU0sIilDBcLLVVperDgalwDnGFjBz5FvhkIIuBQnR
TChtwLCaoNoys/7Z7XeCNpbomcD6aM1zuRV45jSti7Rjfk3IY4TNe6FAAldk2q8q
r7zOtLyCdcFZfCL/lkNcOrLwDlNr7De7+fwz/u9h2kUkw1pUPWzuyxWWooqvWl6b
AqNxkK/fhFQ91DSWRexnQL3lXUoeMddvuldIfbLW1pA/UnmExcESPGl8mTlG4ui/
imckL8w96QbIxrdi4K6i80Mu6utnvAEAf+m0P3eOJgnUzrstbYDls9tXrH2pfFNy
VYcSM+JsRK4RST8Ey67o2aQMYlIWLuAHf/vjxM/DVrgp2cF/d0s03RbQKnDn0QuG
mBd0twDvryQLShnt/tvXW0iN+S3jAYB79oCENj5EX5LNRRVWnox7DoUuki8fodCT
VhtK26xUcT+DaI75ZSbmRy66jzjNhD+dnI7QF+YXZ90cuZMEhzrTjbDs3IVdSThu
ybUnDgHsac6HH2Qrds2b/OElKqJq4p0HrYXMTWLvRXkRUpT3U4D8E7RvssnkU/tB
RK5SOuW2EslufQV2KNZEwHfofbJRtiPZyTBBlwmyARHeGxCNvgHE1QAzLo7rkLGH
Ox9mrquQyPrz8TVBwbBoNt+DOO8G1AfJVQkEDyP9JmGVjrHC/H2pNsois2W+dHRt
pTVZ3sYf81s/Zi+SKwxhUIEy7dZ/E4+Dsstw+cWLhu5YHnGXOrYOt4aBP88WblJL
DzV/ysbXIe9Z2JK0qMCeYphkgLIctjVJtT8D6TEpq3xTm8mQmbEbPRK1w4J8Towy
GaMYac/r9an6SDbikNCvSHBQm33TIr1g/BGpvWr3gwk336ZNco6XKf5iQhk3V7zp
3azlCgd7d7r0lxH4nyENKzKGxl6gkJB3/U4/a8kl6P/hY1yv19oFFyiGupTcsyI6
mgHHPxYaGp5DEX9wroUIifXQHoVHRNrRllQw4o7QxWtrWCS3+7tElcjwg1Q6hxyc
RbrEgMRZNF2AWvyiRN4yuy+wUdHbWQzKaw8XdL6S7WxHeeGj9nyAMUesr0616ajX
JYuYkmYh4G6NJKopTflMty6CbeTqA6PaWdEfXL3lGLRRFCNx0idVhjPfXrw9fU7A
`pragma protect end_protected
