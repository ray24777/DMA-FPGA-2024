//////////////////////////////////////////////////////////////
//  Copyright(c) 2011-2022 Anlogic, Inc.
//  All Right Reserved.
//////////////////////////////////////////////////////////////
//  Company       : Anlogic
//  Filename      : pcie_support.v
//  Author        : Dexin - dexin.guo@anlogic.com
//  Last Modified : 2023-07-26 11:12:21
//  Create        : 2023-06-16 14:58:25
//  Description   :
//
///////////////////////////////////////////////////////////////

`timescale 1ns/1ns


`ifdef DEBUG_MODE
	`include "para_def.vh"
`endif
module pcie_support(

    input   wire                refclk_p                        ,
    input   wire                refclk_n                        ,
    output  wire    [3:0]       txp                             ,
    output  wire    [3:0]       txn                             ,
    input   wire    [3:0]       rxp                             ,
    input   wire    [3:0]       rxn                             ,

    // client0 user interface

    input   wire    [127:0]     client0_tlp_data                ,
    input   wire    [63:0]      client0_tlp_addr                ,
    input   wire    [15:0]      client0_remote_req_id           ,
    input   wire    [7:0]       client0_tlp_byte_en             ,
    input   wire    [11:0]      client0_cpl_byte_cnt            ,
    input   wire                client0_addr_align_en           ,
    input   wire    [2:0]       client0_tlp_tc                  ,
    input   wire    [2:0]       client0_tlp_attr                ,
    input   wire    [2:0]       client0_cpl_status              ,
    input   wire                client0_cpl_bcm                 ,
    input   wire                client0_tlp_dv                  ,
    input   wire                client0_tlp_eot                 ,
    input   wire                client0_tlp_bad_eot             ,
    input   wire                client0_tlp_hv                  ,
    input   wire    [4:0]       client0_tlp_type                ,
    input   wire    [1:0]       client0_tlp_fmt                 ,
    input   wire                client0_tlp_td                  ,
    input   wire    [12:0]      client0_tlp_byte_len            ,
    input   wire    [9:0]       client0_tlp_tid                 ,
    input   wire                client0_tlp_ep                  ,
    input   wire                client0_tlp_func_num            ,
    input   wire    [1:0]       client0_tlp_vfunc_num           ,
    input   wire    [1:0]       client0_tlp_ats                 ,
    input   wire    [7:0]       client0_tlp_st                  ,
    input   wire                client0_tlp_vfunc_active        ,
    input   wire                client0_tlp_nw                  ,
    input   wire                client0_tlp_th                  ,
    input   wire    [1:0]       client0_tlp_ph                  ,
    input   wire                client0_tlp_atu_bypass          ,
    input   wire    [9:0]       client0_cpl_lookup_id           ,
    output  wire                xadm_client0_halt               ,

    // client1 user interface

    input   wire    [127:0]     client1_tlp_data                ,
    input   wire    [63:0]      client1_tlp_addr                ,
    input   wire    [15:0]      client1_remote_req_id           ,
    input   wire    [7:0]       client1_tlp_byte_en             ,
    input   wire    [11:0]      client1_cpl_byte_cnt            ,
    input   wire                client1_addr_align_en           ,
    input   wire    [2:0]       client1_tlp_tc                  ,
    input   wire    [2:0]       client1_tlp_attr                ,
    input   wire    [2:0]       client1_cpl_status              ,
    input   wire                client1_cpl_bcm                 ,
    input   wire                client1_tlp_dv                  ,
    input   wire                client1_tlp_eot                 ,
    input   wire                client1_tlp_bad_eot             ,
    input   wire                client1_tlp_hv                  ,
    input   wire    [4:0]       client1_tlp_type                ,
    input   wire    [1:0]       client1_tlp_fmt                 ,
    input   wire                client1_tlp_td                  ,
    input   wire    [12:0]      client1_tlp_byte_len            ,
    input   wire    [9:0]       client1_tlp_tid                 ,
    input   wire                client1_tlp_ep                  ,
    input   wire                client1_tlp_func_num            ,
    input   wire    [1:0]       client1_tlp_vfunc_num           ,
    input   wire    [1:0]       client1_tlp_ats                 ,
    input   wire    [7:0]       client1_tlp_st                  ,
    input   wire                client1_tlp_vfunc_active        ,
    input   wire                client1_tlp_nw                  ,
    input   wire                client1_tlp_th                  ,
    input   wire    [1:0]       client1_tlp_ph                  ,
    input   wire                client1_tlp_atu_bypass          ,
    input   wire    [9:0]       client1_cpl_lookup_id           ,
    output  wire                xadm_client1_halt               ,
    // trgt user interface
    output  wire                radm_trgt1_dv                   ,
    output  wire                radm_trgt1_hv                   ,
    output  wire                radm_trgt1_eot                  ,
    output  wire                radm_trgt1_tlp_abort            ,
    output  wire                radm_trgt1_dllp_abort           ,
    output  wire                radm_trgt1_ecrc_err             ,
    output  wire    [3:0]       radm_trgt1_dwen                 ,
    output  wire    [1:0]       radm_trgt1_fmt                  ,
    output  wire    [2:0]       radm_trgt1_attr                 ,
    output  wire                radm_trgt1_func_num             ,
    output  wire    [4:0]       radm_trgt1_type                 ,
    output  wire    [2:0]       radm_trgt1_tc                   ,
    output  wire    [15:0]      radm_trgt1_reqid                ,
    output  wire    [127:0]     radm_trgt1_data                 ,
    output  wire    [3:0]       radm_trgt1_first_be             ,
    output  wire    [3:0]       radm_trgt1_last_be              ,
    output  wire    [63:0]      radm_trgt1_addr                 ,
    output  wire    [1:0]       radm_trgt1_vfunc_num            ,
    output  wire                radm_trgt1_vfunc_active         ,
    output  wire                radm_trgt1_td                   ,
    output  wire                radm_trgt1_poisoned             ,
    output  wire                radm_trgt1_hdr_uppr_bytes_valid ,
    output  wire                radm_trgt1_rom_in_range         ,
    output  wire                radm_trgt1_io_req_in_range      ,
    output  wire    [63:0]      radm_trgt1_hdr_uppr_bytes       ,
    output  wire    [2:0]       radm_trgt1_in_membar_range      ,
    output  wire    [2:0]       radm_trgt1_cpl_status           ,
    output  wire    [1:0]       radm_trgt1_ats                  ,
    output  wire    [9:0]       radm_trgt1_tag                  ,
    output  wire    [9:0]       radm_trgt1_dw_len               ,
    output  wire                radm_trgt1_nw                   ,
    output  wire                radm_trgt1_th                   ,
    output  wire    [1:0]       radm_trgt1_ph                   ,
    output  wire    [7:0]       radm_trgt1_st                   ,
    output  wire    [11:0]      radm_trgt1_byte_cnt             ,
    output  wire                radm_trgt1_bcm                  ,
    output  wire    [2:0]       radm_trgt1_vc                   ,
    output  wire    [15:0]      radm_trgt1_cmpltr_id            ,
    output  wire                radm_trgt1_cpl_last             ,
    output  wire    [2:0]       radm_grant_tlp_type             ,
    output  wire    [1:0]       radm_trgt1_atu_sloc_match       ,
    output  wire    [1:0]       radm_trgt1_atu_cbuf_err         ,
    output  wire    [9:0]       trgt_lookup_id                  ,
    output  wire                trgt_lookup_empty               ,
    input   wire                trgt1_radm_halt                 ,
    input   wire    [2:0]       trgt1_radm_pkt_halt             ,
    
    // radm_bypass user interface
    output  wire    [127:0]     radm_bypass_data                ,
    output  wire    [3:0]       radm_bypass_dwen                ,
    output  wire                radm_bypass_dv                  ,
    output  wire                radm_bypass_hv                  ,
    output  wire                radm_bypass_eot                 ,
    output  wire                radm_bypass_dllp_abort          ,
    output  wire                radm_bypass_tlp_abort           ,
    output  wire                radm_bypass_ecrc_err            ,
    output  wire    [63:0]      radm_bypass_addr                ,
    output  wire    [1:0]       radm_bypass_fmt                 ,
    output  wire    [2:0]       radm_bypass_tc                  ,
    output  wire    [2:0]       radm_bypass_attr                ,
    output  wire    [15:0]      radm_bypass_reqid               ,
    output  wire    [4:0]       radm_bypass_type                ,
    output  wire    [9:0]       radm_bypass_tag                 ,
    output  wire                radm_bypass_func_num            ,
    output  wire    [1:0]       radm_bypass_vfunc_num           ,
    output  wire                radm_bypass_vfunc_active        ,
    output  wire                radm_bypass_td                  ,
    output  wire                radm_bypass_poisoned            ,
    output  wire    [9:0]       radm_bypass_dw_len              ,
    output  wire                radm_bypass_rom_in_range        ,
    output  wire    [3:0]       radm_bypass_first_be            ,
    output  wire    [3:0]       radm_bypass_last_be             ,
    output  wire                radm_bypass_io_req_in_range     ,
    output  wire    [2:0]       radm_bypass_in_membar_range     ,
    output  wire                radm_bypass_cpl_last            ,
    output  wire    [2:0]       radm_bypass_cpl_status          ,
    output  wire    [7:0]       radm_bypass_st                  ,
    output  wire    [15:0]      radm_bypass_cmpltr_id           ,
    output  wire    [11:0]      radm_bypass_byte_cnt            ,
    output  wire    [1:0]       radm_bypass_ats                 ,
    output  wire                radm_bypass_th                  ,
    output  wire    [1:0]       radm_bypass_ph                  ,
    output  wire                radm_bypass_bcm                 ,

    // elbi user interface
    output  wire    [31:0]      lbc_ext_addr                    ,
    output  wire    [1:0]       lbc_ext_cs                      ,
    output  wire    [3:0]       lbc_ext_wr                      ,
    output  wire                lbc_ext_rom_access              ,
    output  wire                lbc_ext_io_access               ,
    output  wire    [31:0]      lbc_ext_dout                    ,
    output  wire    [2:0]       lbc_ext_bar_num                 ,
    output  wire                lbc_ext_vfunc_active            ,
    output  wire    [1:0]       lbc_ext_vfunc_num               ,
    input   wire    [63:0]      ext_lbc_din                     ,
    input   wire    [1:0]       ext_lbc_ack                     ,

    // ext drp interface
    input   wire    [31:0]      ext_drp_dbi_din                 ,
    input   wire    [3:0]       ext_drp_dbi_wr                  ,
    input   wire    [31:0]      ext_drp_dbi_addr                ,
    input   wire                ext_drp_dbi_cs                  ,
    input   wire                ext_drp_dbi_cs2_exp             ,
    input   wire    [1:0]       ext_drp_dbi_vfunc_num           ,
    input   wire                ext_drp_dbi_vfunc_active        ,
    input   wire    [2:0]       ext_drp_dbi_bar_num             ,
    input   wire                ext_drp_dbi_rom_access          ,
    input   wire                ext_drp_dbi_io_access           ,
    input   wire                ext_drp_dbi_func_num            ,
    input   wire                ext_drp_app_dbi_ro_wr_disable   ,
    output  wire    [31:0]      ext_drp_lbc_dbi_dout            ,
    output  wire                ext_drp_lbc_dbi_ack             ,

    // msi interface
    output  wire                ven_msi_grant                   ,
    input   wire                ven_msi_req                     ,
    input   wire                ven_msi_func_num                ,
    input   wire    [63:0]      cfg_msi_pending                 ,
    input   wire    [1:0]       ven_msi_vfunc_num               ,
    input   wire                ven_msi_vfunc_active            ,
    input   wire    [2:0]       ven_msi_tc                      ,
    input   wire    [4:0]       ven_msi_vector                  ,
    output  wire    [1:0]       cfg_msi_en                      ,
    output  wire    [63:0]      cfg_msi_mask                    ,

    // system interface
    input   wire                app_power_up_rst_n              ,
    input   wire                app_auxclk                      ,
    output  wire                user_clk                        ,
    output  wire                core_clk                        ,
    output  wire                user_link                       ,
    output  wire                rdlh_link_up

);

// ====================================================================
// Parameter/wire/reg
// ====================================================================

    wire                app_perst_n             =1'b1   ;
    wire                app_button_rst_n        =1'b1   ;

    wire    [5:0]       smlh_ltssm_state                ;//synthesis keep

         

// ====================================================================
// Main Code
// ====================================================================


 


//assign drp_dbi_din_core = drp_dbi_din_user;
//assign drp_dbi_wr_core  = drp_dbi_wr_user;
//assign drp_dbi_addr_core = drp_dbi_addr_user;
//assign drp_dbi_cs_core = drp_dbi_cs_user;
//assign drp_dbi_cs2_exp_core = drp_dbi_cs2_exp_user;
//assign drp_dbi_vfunc_num_core = drp_dbi_vfunc_num_user;
//assign drp_dbi_vfunc_active_core = drp_dbi_vfunc_active_user;
//assign drp_dbi_bar_num_core = drp_dbi_bar_num_user;
//assign drp_dbi_rom_access_core = drp_dbi_rom_access_user;
//assign drp_dbi_io_access_core = drp_dbi_io_access_user;
//assign drp_dbi_func_num_core = drp_dbi_func_num_user;
//assign drp_app_dbi_ro_wr_disable_core = drp_app_dbi_ro_wr_disable_user;
//assign drp_lbc_dbi_ack_user = drp_lbc_dbi_ack_core;
//assign drp_lbc_dbi_dout_user = drp_lbc_dbi_dout_core;


//assign lbc_ext_addr = lbc_ext_addr_core;
//assign lbc_ext_cs = lbc_ext_cs_core;
//assign lbc_ext_wr = lbc_ext_wr_core;
//assign lbc_ext_rom_access = lbc_ext_rom_access_core;
//assign lbc_ext_io_access =  lbc_ext_io_access_core;
//assign lbc_ext_dout =  lbc_ext_dout_core;
//assign lbc_ext_bar_num = lbc_ext_bar_num_core;
//assign lbc_ext_vfunc_active = lbc_ext_vfunc_active_core;
//assign lbc_ext_vfunc_num = lbc_ext_vfunc_num_core;
//assign ext_lbc_din_core = ext_lbc_din;
//assign ext_lbc_ack_core = ext_lbc_ack;

//--------------------------------------------
// pcie ip inst
//--------------------------------------------  

pcie_ep_core
#(
        .SIM_MODE(0)
) 
u_pcie_ep_core 
(
        .refclk_p                          (refclk_p                          ),
        .refclk_n                          (refclk_n                          ),
        .txp                               (txp                               ),
        .txn                               (txn                               ),
        .rxp                               (rxp                               ),
        .rxn                               (rxn                               ),
        .client0_tlp_data                  (client0_tlp_data                  ),
        .client0_tlp_addr                  (client0_tlp_addr                  ),
        .client0_remote_req_id             (client0_remote_req_id             ),
        .client0_tlp_byte_en               (client0_tlp_byte_en               ),
        .client0_cpl_byte_cnt              (client0_cpl_byte_cnt              ),
        .client0_addr_align_en             (client0_addr_align_en             ),
        .client0_tlp_tc                    (client0_tlp_tc                    ),
        .client0_tlp_attr                  (client0_tlp_attr                  ),
        .client0_cpl_status                (client0_cpl_status                ),
        .client0_cpl_bcm                   (client0_cpl_bcm                   ),
        .client0_tlp_dv                    (client0_tlp_dv                    ),
        .client0_tlp_eot                   (client0_tlp_eot                   ),
        .client0_tlp_bad_eot               (client0_tlp_bad_eot               ),
        .client0_tlp_hv                    (client0_tlp_hv                    ),
        .client0_tlp_type                  (client0_tlp_type                  ),
        .client0_tlp_fmt                   (client0_tlp_fmt                   ),
        .client0_tlp_td                    (client0_tlp_td                    ),
        .client0_tlp_byte_len              (client0_tlp_byte_len              ),
        .client0_tlp_tid                   (client0_tlp_tid                   ),
        .client0_tlp_ep                    (client0_tlp_ep                    ),
        .client0_tlp_func_num              (client0_tlp_func_num              ),
        .client0_tlp_vfunc_num             (client0_tlp_vfunc_num             ),
        .client0_tlp_ats                   (client0_tlp_ats                   ),
        .client0_tlp_st                    (client0_tlp_st                    ),
        .client0_tlp_vfunc_active          (client0_tlp_vfunc_active          ),
        .client0_tlp_nw                    (client0_tlp_nw                    ),
        .client0_tlp_th                    (client0_tlp_th                    ),
        .client0_tlp_ph                    (client0_tlp_ph                    ),
        .client0_tlp_atu_bypass            (client0_tlp_atu_bypass            ),
        .client1_tlp_data                  (client1_tlp_data                  ),
        .client1_tlp_addr                  (client1_tlp_addr             ),
        .client1_remote_req_id             (client1_remote_req_id        ),
        .client1_tlp_byte_en               (client1_tlp_byte_en          ),
        .client1_cpl_byte_cnt              (client1_cpl_byte_cnt         ),
        .client1_addr_align_en             (client1_addr_align_en        ),
        .client1_tlp_tc                    (client1_tlp_tc               ),
        .client1_tlp_attr                  (client1_tlp_attr             ),
        .client1_cpl_status                (client1_cpl_status           ),
        .client1_cpl_bcm                   (client1_cpl_bcm              ),
        .client1_tlp_dv                    (client1_tlp_dv               ),
        .client1_tlp_eot                   (client1_tlp_eot              ),
        .client1_tlp_bad_eot               (client1_tlp_bad_eot          ),
        .client1_tlp_hv                    (client1_tlp_hv               ),
        .client1_tlp_type                  (client1_tlp_type             ),
        .client1_tlp_fmt                   (client1_tlp_fmt              ),
        .client1_tlp_td                    (client1_tlp_td               ),
        .client1_tlp_byte_len              (client1_tlp_byte_len         ),
        .client1_tlp_tid                   (client1_tlp_tid              ),
        .client1_tlp_ep                    (client1_tlp_ep               ),
        .client1_tlp_func_num              (client1_tlp_func_num         ),
        .client1_tlp_vfunc_num             (client1_tlp_vfunc_num        ),
        .client1_tlp_ats                   (client1_tlp_ats              ),
        .client1_tlp_st                    (client1_tlp_st               ),
        .client1_tlp_vfunc_active          (client1_tlp_vfunc_active     ),
        .client1_tlp_nw                    (client1_tlp_nw               ),
        .client1_tlp_th                    (client1_tlp_th               ),
        .client1_tlp_ph                    (client1_tlp_ph               ),
        .client1_tlp_atu_bypass            (client1_tlp_atu_bypass       ),
        .ext_lbc_din                       (ext_lbc_din                  ),
        .ext_lbc_ack                       (ext_lbc_ack                  ),
        .sys_atten_button_pressed          (2'b0                              ),
        .sys_pre_det_state                 (2'b0                              ),
        .sys_mrl_sensor_state              (2'b0                              ),
        .sys_pwr_fault_det                 (2'b0                              ),
        .sys_mrl_sensor_chged              (2'b0                              ),
        .sys_pre_det_chged                 (2'b0                              ),
        .sys_cmd_cpled_int                 (2'b0                              ),
        .sys_eml_interlock_engaged         (2'b0                              ),
        .rx_lane_flip_en                   (1'b0                              ),
        .tx_lane_flip_en                   (1'b0                              ),
        .app_req_retry_en                  (1'b0                              ),
        .app_sris_mode                     (1'b1                              ),
        .app_vf_req_retry_en               (4'b0                              ),
        .app_pf_req_retry_en               (2'b0                              ),
        .app_unlock_msg                    (1'b0                              ),
        .app_hdr_log                       (128'b0                            ),
        .app_err_bus                       (13'b0                             ),
        .app_err_advisory                  (1'b0                              ),
        .app_err_func_num                  (1'b0                              ),
        .app_err_vfunc_active              (1'b0                              ),
        .app_hdr_valid                     (1'b0                              ),
        .app_err_vfunc_num                 (2'b0                              ),
        .client0_cpl_lookup_id             (client0_cpl_lookup_id             ),
        .client1_cpl_lookup_id             (client1_cpl_lookup_id             ),
        .app_perst_n                       (app_perst_n                       ),
        .app_power_up_rst_n                (app_power_up_rst_n                ),
        .app_button_rst_n                  (app_button_rst_n                  ),
        //.app_app_ltssm_enable              (app_app_ltssm_enable              ),
        .app_auxclk                        (app_auxclk                        ),
        .drp_dbi_din                       (ext_drp_dbi_din                  ),
        .drp_dbi_wr                        (ext_drp_dbi_wr                   ),
        .drp_dbi_addr                      (ext_drp_dbi_addr                 ),
        .drp_dbi_cs                        (ext_drp_dbi_cs                   ),
        .drp_dbi_cs2_exp                   (ext_drp_dbi_cs2_exp              ),
        .drp_dbi_vfunc_num                 (ext_drp_dbi_vfunc_num            ),
        .drp_dbi_vfunc_active              (ext_drp_dbi_vfunc_active         ),
        .drp_dbi_bar_num                   (ext_drp_dbi_bar_num              ),
        .drp_dbi_rom_access                (ext_drp_dbi_rom_access           ),
        .drp_dbi_io_access                 (ext_drp_dbi_io_access            ),
        .drp_dbi_func_num                  (ext_drp_dbi_func_num             ),
        .drp_app_dbi_ro_wr_disable         (ext_drp_app_dbi_ro_wr_disable    ),
        .phy_cr_para_clk                   (app_auxclk                        ),
        .xadm_client0_halt                 (xadm_client0_halt            ),
        .xadm_client1_halt                 (xadm_client1_halt            ),
        .radm_bypass_data                  (radm_bypass_data             ),
        .radm_bypass_dwen                  (radm_bypass_dwen             ),
        .radm_bypass_dv                    (radm_bypass_dv               ),
        .radm_bypass_hv                    (radm_bypass_hv               ),
        .radm_bypass_eot                   (radm_bypass_eot              ),
        .radm_bypass_dllp_abort            (radm_bypass_dllp_abort       ),
        .radm_bypass_tlp_abort             (radm_bypass_tlp_abort        ),
        .radm_bypass_ecrc_err              (radm_bypass_ecrc_err         ),
        .radm_bypass_addr                  (radm_bypass_addr             ),
        .radm_bypass_fmt                   (radm_bypass_fmt              ),
        .radm_bypass_tc                    (radm_bypass_tc               ),
        .radm_bypass_attr                  (radm_bypass_attr             ),
        .radm_bypass_reqid                 (radm_bypass_reqid            ),
        .radm_bypass_type                  (radm_bypass_type             ),
        .radm_bypass_tag                   (radm_bypass_tag              ),
        .radm_bypass_func_num              (radm_bypass_func_num         ),
        .radm_bypass_vfunc_num             (radm_bypass_vfunc_num        ),
        .radm_bypass_vfunc_active          (radm_bypass_vfunc_active     ),
        .radm_bypass_td                    (radm_bypass_td               ),
        .radm_bypass_poisoned              (radm_bypass_poisoned         ),
        .radm_bypass_dw_len                (radm_bypass_dw_len           ),
        .radm_bypass_rom_in_range          (radm_bypass_rom_in_range     ),
        .radm_bypass_first_be              (radm_bypass_first_be         ),
        .radm_bypass_last_be               (radm_bypass_last_be          ),
        .radm_bypass_io_req_in_range       (radm_bypass_io_req_in_range  ),
        .radm_bypass_in_membar_range       (radm_bypass_in_membar_range  ),
        .radm_bypass_cpl_last              (radm_bypass_cpl_last         ),
        .radm_bypass_cpl_status            (radm_bypass_cpl_status       ),
        .radm_bypass_st                    (radm_bypass_st               ),
        .radm_bypass_cmpltr_id             (radm_bypass_cmpltr_id        ),
        .radm_bypass_byte_cnt              (radm_bypass_byte_cnt         ),
        .radm_bypass_ats                   (radm_bypass_ats              ),
        .radm_bypass_th                    (radm_bypass_th               ),
        .radm_bypass_ph                    (radm_bypass_ph               ),
        .radm_bypass_bcm                   (radm_bypass_bcm              ),
//        .radm_trgt1_dv                     (radm_trgt1_dv                ),
//        .radm_trgt1_hv                     (radm_trgt1_hv                ),
//        .radm_trgt1_eot                    (radm_trgt1_eot               ),
//        .radm_trgt1_tlp_abort              (radm_trgt1_tlp_abort         ),
//        .radm_trgt1_dllp_abort             (radm_trgt1_dllp_abort        ),
//        .radm_trgt1_ecrc_err               (radm_trgt1_ecrc_err          ),
//        .radm_trgt1_dwen                   (radm_trgt1_dwen              ),
//        .radm_trgt1_fmt                    (radm_trgt1_fmt               ),
//        .radm_trgt1_attr                   (radm_trgt1_attr              ),
//        .radm_trgt1_func_num               (radm_trgt1_func_num          ),
//        .radm_trgt1_type                   (radm_trgt1_type              ),
//        .radm_trgt1_tc                     (radm_trgt1_tc                ),
//        .radm_trgt1_reqid                  (radm_trgt1_reqid             ),
//        .radm_trgt1_data                   (radm_trgt1_data              ),
//        .radm_trgt1_first_be               (radm_trgt1_first_be          ),
//        .radm_trgt1_last_be                (radm_trgt1_last_be           ),
//        .radm_trgt1_addr                   (radm_trgt1_addr              ),
//        .radm_trgt1_vfunc_num              (radm_trgt1_vfunc_num         ),
//        .radm_trgt1_vfunc_active           (radm_trgt1_vfunc_active      ),
//        .radm_trgt1_td                     (radm_trgt1_td                ),
//        .radm_trgt1_poisoned               (radm_trgt1_poisoned          ),
//        .radm_trgt1_hdr_uppr_bytes_valid   (radm_trgt1_hdr_uppr_bytes_valid),
//        .radm_trgt1_rom_in_range           (radm_trgt1_rom_in_range      ),
//        .radm_trgt1_io_req_in_range        (radm_trgt1_io_req_in_range   ),
//        .radm_trgt1_hdr_uppr_bytes         (radm_trgt1_hdr_uppr_bytes    ),
//        .radm_trgt1_in_membar_range        (radm_trgt1_in_membar_range   ),
//        .radm_trgt1_cpl_status             (radm_trgt1_cpl_status        ),
//        .radm_trgt1_ats                    (radm_trgt1_ats               ),
//        .radm_trgt1_tag                    (radm_trgt1_tag               ),
//        .radm_trgt1_dw_len                 (radm_trgt1_dw_len            ),
//        .radm_trgt1_nw                     (radm_trgt1_nw                ),
//        .radm_trgt1_th                     (radm_trgt1_th                ),
//        .radm_trgt1_ph                     (radm_trgt1_ph                ),
//        .radm_trgt1_st                     (radm_trgt1_st                ),
//        .radm_trgt1_byte_cnt               (radm_trgt1_byte_cnt          ),
//        .radm_trgt1_bcm                    (radm_trgt1_bcm               ),
//        .radm_trgt1_vc                     (radm_trgt1_vc                ),
//        .radm_trgt1_cmpltr_id              (radm_trgt1_cmpltr_id         ),
//        .radm_trgt1_cpl_last               (radm_trgt1_cpl_last          ),
//        .radm_grant_tlp_type               (radm_grant_tlp_type          ),
//        .radm_trgt1_atu_sloc_match         (radm_trgt1_atu_sloc_match    ),
//        .radm_trgt1_atu_cbuf_err           (radm_trgt1_atu_cbuf_err      ),
        .training_rst_n                    (),
        .lbc_ext_addr                      (lbc_ext_addr                 ),
        .lbc_ext_cs                        (lbc_ext_cs                   ),
        .lbc_ext_wr                        (lbc_ext_wr                   ),
        .lbc_ext_rom_access                (lbc_ext_rom_access           ),
        .lbc_ext_io_access                 (lbc_ext_io_access            ),
        .lbc_ext_dout                      (lbc_ext_dout                 ),
        .lbc_ext_bar_num                   (lbc_ext_bar_num              ),
        .lbc_ext_vfunc_active              (lbc_ext_vfunc_active         ),
        .lbc_ext_vfunc_num                 (lbc_ext_vfunc_num            ),
        .rdlh_link_up                      (rdlh_link_up                      ),
        .cfg_vf_bme                        (),
        .radm_vendor_msg                   (),
        .radm_msg_payload                  (),
        .radm_msg_req_id                   (),
        .cfg_send_cor_err                  (),
        .cfg_send_nf_err                   (),
        .cfg_send_f_err                    (),
        .cfg_link_eq_req_int               (),
        .smlh_req_rst_not                  (),
        .link_req_rst_not                  (),
        .radm_msg_unlock                   (),
        .smlh_ltssm_state                  (smlh_ltssm_state                  ),
        .radm_cpl_timeout                  (),
        .radm_timeout_func_num             (),
        .radm_timeout_vfunc_num            (),
        .radm_timeout_vfunc_active         (),
        .radm_timeout_cpl_tc               (),
        .radm_timeout_cpl_attr             (),
        .radm_timeout_cpl_tag              (),
        .radm_timeout_cpl_len              (),
        .pm_xtlh_block_tlp                 (),
        .cfg_phy_control                   (),
        .cfg_hw_auto_sp_dis                (),
        .smlh_ltssm_state_rcvry_eq         (),
        .trgt_cpl_timeout                  (),
        .trgt_timeout_cpl_func_num         (),
        .trgt_timeout_cpl_vfunc_num        (),
        .trgt_timeout_cpl_vfunc_active     (),
        .trgt_timeout_cpl_tc               (),
        .trgt_timeout_cpl_attr             (),
        .trgt_timeout_cpl_len              (),
        .trgt_timeout_lookup_id            (),
        .trgt_lookup_id                    (trgt_lookup_id                    ),
        .trgt_lookup_empty                 (trgt_lookup_empty                 ),
        .cfg_reg_serren                    (),
        .cfg_cor_err_rpt_en                (),
        .cfg_nf_err_rpt_en                 (),
        .cfg_f_err_rpt_en                  (),
        .cfg_uncor_internal_err_sts        (),
        .cfg_rcvr_overflow_err_sts         (),
        .cfg_fc_protocol_err_sts           (),
        .cfg_mlf_tlp_err_sts               (),
        .cfg_surprise_down_er_sts          (),
        .cfg_dl_protocol_err_sts           (),
        .cfg_ecrc_err_sts                  (),
        .cfg_corrected_internal_err_sts    (),
        .cfg_replay_number_rollover_err_sts(),
        .cfg_replay_timer_timeout_err_sts  (),
        .cfg_bad_dllp_err_sts              (),
        .cfg_bad_tlp_err_sts               (),
        .cfg_rcvr_err_sts                  (),
        .ven_msi_grant                     (ven_msi_grant                     ),
        .ven_msi_req                       (ven_msi_req                       ),
        .ven_msi_func_num                  (ven_msi_func_num                  ),
        .cfg_msi_pending                   (cfg_msi_pending                   ),
        .ven_msi_vfunc_num                 (ven_msi_vfunc_num                 ),
        .ven_msi_vfunc_active              (ven_msi_vfunc_active              ),
        .ven_msi_tc                        (ven_msi_tc                        ),
        .ven_msi_vector                    (ven_msi_vector                    ),
        .cfg_msi_en                        (cfg_msi_en                        ),
        .cfg_msi_mask                      (cfg_msi_mask                      ),
        .core_rst_n                        (core_rst_n                        ),
        .drp_lbc_dbi_dout                  (ext_drp_lbc_dbi_dout              ),
        .drp_lbc_dbi_ack                   (ext_drp_lbc_dbi_ack               ),
        .core_clk                          (core_clk                          ),
        .user_link                         (user_link                         ),
        .user_clk                          (user_clk                          ),
        .muxd_aux_clk                      (),
        .muxd_aux_clk_g                    ()

) ;




endmodule
