/*===========================================*\
Filename         : sgdma_ip.v
Project name     : sgdma_subsys_tst
Description      : Merge all submodules of DMA controller core.
Called by        : sgdma_subsys.v
Email            : bingsong.wang@anlogic.com
Modified         : v1.0 Original version,accomplish the basic functions;20210412	  
Copyright(c)Shanghai Anlu Information Technology Co.,Ltd
\*===========================================*/
`ifdef DEBUG_MODE
	`include "../def/para_def.vh"
`else
    `include "../def/para_def.vh"
`endif
module sgdma_ip(
	input   core_rst_n,
	input   core_clk,
	
	input   [1:0]    lbc_ext_cs_i,
    output  [1:0]    ext_lbc_ack_o,
    input   [31:0]   lbc_ext_addr_i,
    input   [3:0]    lbc_ext_wr_i,
    output  [63:0]   ext_lbc_din_o, 
    input   [31:0]   lbc_ext_dout_i,
	input            lbc_ext_rom_access_i,
	input            lbc_ext_io_access_i,
	input   [2:0]    lbc_ext_bar_num_i,
	input            lbc_ext_vfunc_active_i,
	input   [1:0]    lbc_ext_vfunc_num_i,
	
	output   client0_addr_align_en_o,
	output   [`HEADER_WIDTH-1:0] client0_tlp_header_o,
	output   client0_tlp_dv_o,
	output   client0_tlp_eot_o,
	output   client0_tlp_bad_eot_o,
	output   client0_tlp_hv_o,
	output   [12:0]   client0_tlp_byte_len_o,
	output   [`DATA_WIDTH-1:0]   client0_tlp_data_o,
	output   client0_tlp_func_num_o,
	output   [1:0]   client0_tlp_vfunc_num_o,
	output   client0_tlp_vfunc_active_o,
	input    xadm_client0_halt_i,
	output   client0_tlp_atu_bypass_o,
	
	output   client1_addr_align_en_o,
	output   [`HEADER_WIDTH-1:0] client1_tlp_header_o,
	output   client1_tlp_dv_o,
	output   client1_tlp_eot_o,
	output   client1_tlp_bad_eot_o,
	output   client1_tlp_hv_o,
	output   [12:0]   client1_tlp_byte_len_o,
	output   [`DATA_WIDTH-1:0]   client1_tlp_data_o,
	output   client1_tlp_func_num_o,
	output   [1:0]   client1_tlp_vfunc_num_o,
	output   client1_tlp_vfunc_active_o,
	input    xadm_client1_halt_i,
	output   client1_tlp_atu_bypass_o,
	
	input    radm_bypass_dv_i,
	input    radm_bypass_hv_i,
	input    radm_bypass_eot_i,
	input    [`DATA_WIDTH-1:0]     radm_bypass_data_i,
	input    [`HEADER_WIDTH-1:0]   radm_bypass_header_i,//pos&non_pos 4DW,cpl 3DW. 
	input    [1:0]  radm_bypass_dwen_i,
	input    radm_bypass_cpl_last_i,
	input    radm_bypass_dllp_abort_i,
	input    radm_bypass_tlp_abort_i,
	input    radm_bypass_ecrc_err_i,
	input    radm_bypass_func_num_i,
	input    [1:0]  radm_bypass_vfunc_num_i,
	input    radm_bypass_vfunc_active_i,
	input    radm_bypass_io_req_in_range_i,
	input    [2:0]  radm_bypass_in_membar_range_i,
	input    radm_bypass_rom_in_range_i,
`ifdef AXIL_MBUS0_EN	
	output 	[31:0]   m_axil_awaddr_o,
	output 	[2:0]    m_axil_awprot_o,	
	output 	m_axil_awvalid_o,	
	input  	m_axil_awready_i,	
	output 	[31:0]   m_axil_wdata_o,	
	output 	[3:0]    m_axil_wstrb_o,	
	output 	m_axil_wvalid_o,	
	input  	m_axil_wready_i,	
	input  	m_axil_bvalid_i,	
	input  	[1:0] m_axil_bresp_i,	
	output 	m_axil_bready_o,
	output 	[31:0]   m_axil_araddr_o,	
	output 	[2:0]    m_axil_arprot_o,	
	output 	m_axil_arvalid_o,	
	input  	m_axil_arready_i,	
	input  	[31:0]   m_axil_rdata_i,	
	input  	[1:0]    m_axil_rresp_i,	
	input  	m_axil_rvalid_i,		
	output 	m_axil_rready_o,	
`endif	
`ifdef AXIL_SBUS0_EN
	input   [31:0]   s_axil_awaddr_i,
	input   [2:0]    s_axil_awprot_i,
	input            s_axil_awvalid_i,	
	output           s_axil_awready_o,	
	input   [31:0]   s_axil_wdata_i,	
	input   [3:0]    s_axil_wstrb_i,	
	input            s_axil_wvalid_i,	
	output           s_axil_wready_o,	
	output           s_axil_bvalid_o,	
	output  [1:0]    s_axil_bresp_o,	
	input            s_axil_bready_i,	
	input   [31:0]   s_axil_araddr_i,	
	input   [2:0]    s_axil_arprot_i,	
	input            s_axil_arvalid_i,	
	output           s_axil_arready_o,	
	output  [31:0]   s_axil_rdata_o,	
	output  [1:0]    s_axil_rresp_o,	
	output           s_axil_rvalid_o,	
	input            s_axil_rready_i,
`endif

`ifdef AXIS_BUS0_EN
	output   s0_axis_tx_rst_o,
    output   m0_axis_rx_rst_o,
    output   s0_axis_tx_run_o,
    output   m0_axis_rx_run_o,
    
	output   s0_axis_tx_tready_o,
    input    [`DATA_WIDTH-1:0]    s0_axis_tx_tdata_i,
    input    [`KEEP_WIDTH-1:0]    s0_axis_tx_tkeep_i,
    input    [`KEEP_WIDTH-1:0]    s0_axis_tx_tuser_i,
    input    s0_axis_tx_tlast_i,
    input    s0_axis_tx_tvalid_i,	
	input    m0_axis_rx_tready_i,
    output   [`DATA_WIDTH-1:0]    m0_axis_rx_tdata_o,
    output   [`KEEP_WIDTH-1:0]    m0_axis_rx_tkeep_o,
    output   [`KEEP_WIDTH-1:0]    m0_axis_rx_tuser_o,
    output   m0_axis_rx_tlast_o,
    output   m0_axis_rx_tvalid_o,
`endif
`ifdef AXIS_BUS1_EN
	output   s1_axis_tx_tready_o,
    input    [`DATA_WIDTH-1:0]    s1_axis_tx_tdata_i,
    input    [`KEEP_WIDTH-1:0]    s1_axis_tx_tkeep_i,
    input    [`KEEP_WIDTH-1:0]    s1_axis_tx_tuser_i,
    input    s1_axis_tx_tlast_i,
    input    s1_axis_tx_tvalid_i,
	input    m1_axis_rx_tready_i,
    output   [`DATA_WIDTH-1:0]    m1_axis_rx_tdata_o,
    output   [`KEEP_WIDTH-1:0]    m1_axis_rx_tkeep_o,
    output   [`KEEP_WIDTH-1:0]    m1_axis_rx_tuser_o,
    output   m1_axis_rx_tlast_o,
    output   m1_axis_rx_tvalid_o,
`endif
`ifdef AXI4_BUS0_EN
	input   m_axi_arready_i,
	output  [3:0] m_axi_arid_o,
	output  [`DATA_WIDTH-1:0] m_axi_araddr_o,
	//specifies the number of data transfers that occur within each burst.
	output  [7:0] m_axi_arlen_o,
	//specifies the maximum number of data bytes to transfer in each beat. 011-8byte,100-16byte
	output  [2:0] m_axi_arsize_o,
	output  [1:0] m_axi_arburst_o,
	output  [2:0] m_axi_arprot_o,
	output  m_axi_arvalid_o,
	output  m_axi_arlock_o,
	output  [3:0] m_axi_arcache_o,
	
	input   [3:0] m_axi_rid_i,
	input   [`DATA_WIDTH-1:0]m_axi_rdata_i,
	input   [1:0] m_axi_rresp_i,
	input   m_axi_rlast_i,
	input   m_axi_rvalid_i,
	output  m_axi_rready_o,
	
	input   m_axi_awready_i,
	output  [3:0] m_axi_awid_o,
	output  [`DATA_WIDTH-1:0] m_axi_awaddr_o,
	output  [7:0] m_axi_awlen_o,
	output  [2:0] m_axi_awsize_o,
	output  [1:0] m_axi_awburst_o,
	output  [2:0] m_axi_awprot_o,
	output  m_axi_awvalid_o,
	output  m_axi_awlock_o,
	output  [3:0] m_axi_awcache_o,
	output  [`DATA_WIDTH-1:0] m_axi_wdata_o,
	output  [7:0] m_axi_wstrb_o,
	input   m_axi_wready_i,
	output  m_axi_wlast_o,
	output  m_axi_wvalid_o,
	input   [3:0] m_axi_bid_i,
	input   [1:0] m_axi_bresp_i,
	input   m_axi_bvalid_i,
	output  m_axi_bready_o,
`endif	
`ifdef USR_IRQ_EN
	input   ven_msi_grant_i,
	input   [1:0]   cfg_msi_en_i,
	input   [63:0]  cfg_msi_mask_i,	
	output  ven_msi_req_o,
	output  ven_msi_func_num_o,
	output  [1:0]   ven_msi_vfunc_num_o,
	output  ven_msi_vfunc_active_o,
	output  [2:0]   ven_msi_tc_o,
	output  [4:0]   ven_msi_vector_o,
	output  [63:0]  cfg_msi_pending_o,
	/*
	input   [1:0]    cfg_int_disable_i,
	input   [15:0]   cfg_int_pin_i,
	input   assert_inta_grt_i,
	input   assert_intb_grt_i,
	input   assert_intc_grt_i,
	input   assert_intd_grt_i,
	input   deassert_inta_grt_i,
	input   deassert_intb_grt_i,
	input   deassert_intc_grt_i,
	input   deassert_intd_grt_i,
	output  [1:0]   sys_int_o,
	*/
	input   [`DMA_USR_IRQ-1:0]   usr_irq_req_i,
	output  [`DMA_USR_IRQ-1:0]   usr_irq_ack_o,
	output  msi_enable_o,
	output  [2:0]   msi_vector_width_o,
`endif
//  output                                  rdscp0_eot_out,
//    output                                rd0_rden_out,
`ifdef CFG_MGMT_EN 
	//---dbi2cfg interface---
	input   rdlh_link_up_i,
	output  [31:0]  drp_dbi_din_o,
    output  [3:0]   drp_dbi_wr_o,
    output  [31:0]  drp_dbi_addr_o,
    output 	        drp_dbi_cs_o,
	output          drp_dbi_cs2_o,
    input   [31:0]  drp_lbc_dbi_dout_i,//  
    input 	        drp_lbc_dbi_ack_i, //  
    output  [1:0]   drp_dbi_vfunc_num_o,	
    output          drp_dbi_vfunc_active_o,
	output          drp_dbi_func_num_o,
	output          drp_dbi_rom_access_o,
	output          drp_dbi_io_access_o,
	output          drp_app_dbi_ro_wr_disable_o,
	output  [2:0]   drp_dbi_bar_num_o,	
	input   [18:0]  cfg_mgmt_addr_i,
	input   cfg_mgmt_write_i,
	input   [31:0]  cfg_mgmt_write_data_i,
	input   [3:0]   cfg_mgmt_byte_enable_i,	
	input   cfg_mgmt_read_i,	
	output  [31:0]  cfg_mgmt_read_data_o,	
	output  cfg_mgmt_read_write_done_o,
	input   cfg_mgmt_type1_cfg_reg_access_i
`endif
);
//---Start encrypt
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
W5846/gfDd0sZaGay37+ny2Pos9Bdt8tc2hMalxoEb7i/ZYujn9oraLkLw4Wp0V+
NowVE/60Ah59BEDoNa0CTnks5BrBgz15TT1K/VZfOiB7AcXcJzUmW+3Kht+5KG6G
0/eVyS9huVvkz/otIpeVhKBsgymtMSqL0RiVsDmqJvc=
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
Vc2l41zIVcUY16oWLyqjVi4D1kZt4yJ3Q1Ll6/nPm963r7Y+guqG4BATmgVDAate
pk3yhJLWoTFtRADTyCVKAXxoswZdBUlspyM7O9ab/EvDr5bPJv3wQ+w9M3iGRoNu
+TXST9LBlVSKcMp/5WI5nG/b+Zj7oG6xhbSsycTu68Bp5qmQ9rYtziZxxInThmzK
3qCebOm55ZS2R3QgTBFhHfJGqKGsPkbgjzp1wRfLWMlqOgPACzDz6Jgp1QmBqegU
3Xfy4xBl9txj3ypxSnfpIun/ysB0VqcO05OFsee+l6M3pfFlF87qq5opkU0xQz6p
VHLrFaxFwafi4xQgz9mVIw==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
SCZXMLPcmNUcLZXI4+rTCV+MxO1zWoQnffiRAmpKhGvoi0A4vuag3wLd7/tr981v
XxabGQT4GR3C8JbZaWQets/m3+WXbaNXEK3qdHCLflrTmhTakY0VXnMzu+YK/r3F
uRT4RXw3Km0WpmPotxMcNDNngy5xB1zeAFzP0Pw6hmE=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
UTwUPQQ2hVYZvzGjGfBh8MwSvWDCWzroVNJUN2UgH9vY3LVcNrSBuMkRkN37qm87
Ag9MlK5t+JtKZfSXZOKUFhbcwibt03kW9MjOi+kZ0PEnHpTkOz1JW6BAyKTO8mt+
LWMK5iuKcnDpnFuemyNitfCjBhSVNNe1rIvXILPHqpJxc4h6yRJQQ9Fj/QKZ9Wx7
FYHVLezpWzJKiMOxEi2UyGQqBN56tbK3I+IsYoeZAOHjWD14kEpG5LwSq6W/HkKC
fbCwDFjxCU567u2fuiXestfar3y/7oEQ2Z/AbsAoVc8K6LiYc5hn9DI+EkzpTcdt
JIxQmuMvjOdbx6Spldfj9w==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
a5UZBC8cMz42WiX7YTlUQ/BORhGIyrasmJ0OQgOgiYfBGf3eG4XwkNy4dNbLJ7ET
B9ZKyf/fwVqlUoasW/HQ2lITt/NrqDGiZDkLxYOzHBylqxTbfvO8k+4W8QlsbkNE
p83R8Y81mkxa6miw8u7jS0zSFZhkWnrfGJMGcEIV2yQ=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 312592)
`pragma protect data_block
cTZ3bXAyZnlxMmRGVjdIU0HRm23Kvkjg3GkZJ9ExprhUBhEGo5bUuWeLW9WHP3jM
zDzCL/M7jDVnLDARIEZMj8vESj2UCYDoPojdwndJW+SbWTyJT2R5uhESaWeDo9nO
RtkbBq8RaYfcCRc/sj2hyvQ/FtPLn9MWx/lESZ+Yd1kP/lZx3aWa8JwA0pOeAE5o
nk4e2cftGrZgPC6Xnhy32te/5SXkap39WEn2vNgVYLQIcbcEo80gOqpD8b0qEaHh
XLl/mEDSCPXNrIR99VlRZwZ6lDMWUxMqm/+btRqSltEtaE2wdO6tingEuR2VYkur
CFUavnI21Cghr1ctDdiGs8/g4arD2Mr6A8Ux995ibCwn/MQSkMCKyIOupW1od36W
lVDcdKmPUR+raWzBekjxW83zhF0CkyLHKm4R3OeKQsLdelHJWuJ5CvZmUXOvC5qi
DNz8yRI1DBtkKZaP/0rvMDWh4CBZzDMfLGcZ4WHf0XFdtB4zydOxGbjjLE6yKnD2
cjXsOcjkVrq7h4HmWJ8I2Myj+LiVMZ4ypJDjaxkMJuBruoGx/wWIW80e20BHSwSJ
DOc20CejGmgwH7EsYGQnMfe6qO7Cu9aCnGvQzy1lYpeu1qNC0AXqXihLkYepjCXB
Bg7Jj/6vQl/Fzk3Up+g2IwZg1p0u5mSmOG36IYyG5CfF5yITORqPF/MZkdLG1c7Y
cE54Cd748vN7vxZUg2RgaebDgli4PzsAZPBD1fG1w4xWJ/krYfX/YhP//ePHbKVQ
nEu+fywvr0ipHDDM1QfOota15Xw0J3+VZH1siMVV2VT6u/RMbcfWQku3utDWafmu
RxvU8/bKrAUMFwiMe5qlB93SOgNvY0wnSSs2mmRfpnSkwwy8qZZ+E4Mu+OH6iO8p
t+Qd16UJUoB7B0Llk3mfdeTApjXO64RFngux73NfSri/6MUX2jRMK5wSrmKvBje6
AbvrXXmrbavJHUtbUMgJxiq6mhiynl+fjC/bIAParmJOzCTK8BpHdJtW+328W+lp
65+V2d14/hoTvQ89qQOIQcOl5e3pO3+9DhEnlca6gLd9Itg4v2Lma5U0UZloW4e5
Ft/bKXRzGoR/l9YEJWn+jacRpUt006lX1szYr+7n5L6xzgzz0O2mG/d6HxJ39X5R
cmd6cOIx7PKsgztSCX/u6FyYnr6EfFk9YaVkSvFeMwIuscuMh+J+UroekARBmrFk
GfDDwN6QDfXZLM0HKQD10AjQDoqmPh+0ifXqr3iIVtYAnOtE/LQaREm5t7Wns8cI
bOba4y4PyrvXW4K/4ucbMrPL053+1C2g7rvN9MvzjgG/QmYzj4pxVK6I/jgAvQGc
PUy9v8kyzB+4bb2zmOXN7ua3/BMyKf1HrV1AlsIh0hIT5jdKt9hdI+Vjd6tkZHZh
/HBU17pxt8iitDgOHMIdVjVdv03CYRuAe2s+ZNqEiM6/gqVKwz9Q7ZM//N1oT4ys
mVRX813O5S09Qh94RRA0GbNPB65U7HiVhPSWHYFUcLWVBF3FQUW3OQftN4/YCgrx
SyQETl7xQ8ZR980wQ+Ko4OPnOTkkOvWsooNZLAA4hRkuflQdy9chf8gE/oDtvRf7
0t4LlzT3dae+CfvDb1oVRsJg9hR4+IFWKfcZSq9rgfzYNfCAiQn0OEfhBuCqkWev
TNGDcxB710IradcXpTBeAWHvj4lruVMzQQQpMDntMXiX30Yxz2BqrJEO1H9h6bmH
/F5Tf6LFKSxSTv3T6zKzSkDav0viEB7KG27Bo3VP4i6SJbSOKVF1XvKmmUggrHuG
LCKw0YWG0JacgKpIFDucnvQ9qJdnLGJFWZYsiNAAQMZRqnNfU7QNNU9tVIK0i8N2
z7rGtxvERQS1JvetiBFWeLZ0KNxoEU+N6Zx7OAAxg5+webkMyztJxTAa/iqzbOOe
m7e3Q4dGxRmsORKmQRjEWoE1oiMCF2BYwG1lE3nDiR0tFR3GyrYEcNpq69qRDlfJ
Xzd6LziPksLJ8nTu3FR7EvdODGuE1yaGb4nrlDf6dtbrcBGF9XoGHq/YkHuvDplJ
Dn4wIhxnb3Au8oJ4UKeo1udA2TP2oiFDZ1YhTHSgh1cXHkfK8hIAcj8QmNvCNpfc
kXbJ+gHd1w4dMzPBhBHIRbd2YEBzVM+k0K1vhbyAu4rys2Q9XTGerr9W04sDE90v
OWfwJK+JtAY7vHpzyHEEfudgv2csGF9dF2EJNRmaO9YTCq9S/FapK6KoHcszLkeQ
zjRHx3REiBM9Fd5KXV6Oabg/s4Iq9o4Hg4kiOfQEBh8fm93jYCwtEUJmXU8L1mog
hhPXg9gaRQclD/KaK/oPe4TR9K/w1u8IHqL+uPKpz8kX1q123KR1gyHeWlnVNYSF
qEwBZorS0XiCvlC4cr+0ZGIRcpHCLBPcuTCiZpzlRbizHwM8HdLvv3Tla9tt2kUD
LYS82LREkON/UvwzRfp0mu3eKtAnQccgmCn8zCToZDgZR6CqNadcZ6bezEmSaGj+
Ap9E6bmCeKOiko0hcnT7rAAkDEweB4oK295r3toB1OZUxWA/LrxxaAJNep7rYFU/
IfphT1zltPt0ooKiyFszpr+XnyXKAZVuoYr054ColKnd7uZKCwez9bmsxbKG3K0p
Bhl/S9Fz4vWkHDHgks7XwWKxCRU/BuL7rkmzfYRtq2FKKiuhloX0b3o9yCpLkhAB
EWlGJBIohXvqHJMsiA7TMqH/aNnMOTOQOkGqDI+ToiDeghWDzFoC1qjYAHfSxCMT
nxdSSVX/PJGy7+KfGAN492n9xBXbQoFzFCfWBheq2/hq87BLle3RmZZguB2h/JgE
55wgE5zIIM/uj0LYW9nRbipoveV9QXajj74j3gnfBPjw9t1nQnlZ26WQY7JhBA5B
7Bag9gMJUDw0hdjsElLZsX/eiVR2Ft65rCmjVipe/0nswiBTXX5d6lTdDa4ZQBQv
EyL/Atbz2irsrNCOrB2+1bJH6/6J6zVWa7fw7cGMKFcKyWZrHIG+nSBgHSRoHk8q
mORpDL8Fnir1iTA/GdyaxLv+LAbatvSsKETJUKj15Ed6+xsmAGAg2DUWT5STEJAM
mRYWZ5tmmY0NdLnneBb40pxzF1xCX12xWA0BsbtVlsWqnqoqEGIxxqjB+NopQhne
T2WOHZnqf8CBVC4Aim3Xc1sGqeAoHzwwa6OPcHb+nI0va8oZ4Wprb9XPriw+sGX1
HerXvrEqIHBoxy3wGUESV/rSE8C0I8tLvY1s+vV5e49okeQ6Obv/LW46K8jnYvwU
n1CV3p0ZujCa/zCmoq0Sz1wNvSpmkx5J80M9b8diWE2cSciHpSfXczcvBPYxyAt1
szdIMuyxXktxSjO71RnXD8pmQEDsNfdDtzCCXFhTZQ6nUh6kZ2hR/Ia5Bw6o32f1
YjKraIzpLAwX/UiZpqhzk4sU+Z/8ZdvhMDzbxYmoohk+81hi2/cPV1Y3mobV8QF5
TO1SZKPo9AU1GaL0LBWgOBemT5K+g976GgtEM3t0s6WeL0eesVkpt1BHTHP3fu04
oM50FbLnTGhPaOPwnBLkMdMwoNzCX0Dwdhjof3pCwx82kG5MM4SKgQS2EC3/qti9
+Q4u2ju3Bz2xJhwGKCmQbRKxITBBEHnezvs888CibmMnKdvy6AaB119LN4ABT6ql
WxN1cM2OrM6GaWRZ1PEBqxbroPvXeZVRwQJ5MKXthmsdRl6HXq/PoRAatyEiaejx
AHFxMSvbbumggAMSJ7vRgLhxVfd2ST2lfP2cYLb2iMF0atrzNHGqoDnCusX7/NAy
CM2XC8v3voTk2YgpfvwSTmoJ4+3VDf813Qrpqo1OTS7leLFhkkdMymuLQYOewNqM
jg67y+8sDIaQM8Fnofo5Q8WzRhJHFlTQ8dd2qPpGT2MG8rijKmGr/MZQA6WTJtnL
ZtTBHEPkgSKrSoXiQwYb+WS7QheLW1iCU2pB2E9aktqZNSnBuWEmEJqWHavhAaqu
euE2u3JBPy4rMpg8P1CtAQM5vixxqflo/Yk/VqUuqRu/SN0Lal+if96LWIuMEviJ
ZeWaSMPOAfKu5L+vKAALpfS98Tyr9dTCg89qR5b5z7mqNUDkkQjsjR6xewdbEVKb
T0/ap3t6f1bicmHcnpAm/qq3l7/U1yTsxE4r5zeCluqfg3zExiQG38j3Dm8u5c5Y
JvXYObnJksiVn8yRGvoYmYyZw/TKj1uCY1FK5gH6pm7dSYjxA1xstTDze2Ke/djO
zCzuqEV0FYjXgA9RGOlo+BuYqLICzFbqiCtuo8MI9aurnK/Ay2VRsmsA1nQ3OiUz
nC8Oeyrna5FVVT12FR7bQpxrLNarbedlrKOJboqnQsh+PFOqThYtN+3q0Qqv8azg
QMuE/A2dlvNmUkGbqnPC9peFrSmsf2j8Y0CloM6BqSEwp8L+xNAe21iue5LM1ZPl
p7NcIyBn/4jPuvKnTJpIIJD9dlxc2OpPbT7gYL85rpmmis8C+gBntZqG5fCSqXOP
ZfXJFstfH/dn/kJkBp+NiMx+V0Ag5nNBAdqcXd/oedeUdISuqK92mnfjHxXQsmcx
+Z+RPuy/OAjdYxz4Q3BW+1Trh0Uc+0oyGuNiYG8YyFSmSzpGVy/StSc2Vn287MSE
oloMEw/tWsguuhp7yaOeKmEKA3I1znztvfSZhzAbcC/b8r2QnPVC69uQBhDogvzA
WPXOWmin8oaVpnUL7UwRVxKddU825hgH8VSvbitTnSxEvtSyHHVFtIZt7rzmDZLz
XgcFLLRnW2W7hHFPPkoEvFjIqRUEHRWGYg5MN1wh794PBPKAO4/NCokGssKjQUL6
Ua/IKOjx4bHCsy+V44O+IYIKCWcnnXcBoylTA3Upro3OOJE+a63qCbVBtXfp5iI2
VnEhdjKfGa+gG8mJVNV3zrCbqamg/szDO6l1wdf+f8+lgHmCBJ1EoJzKzAaZEeYN
zfYA7dTIkn9uQYugTfpnOVHThj5ny0Diilu4u+9vEliN30cdB1Z46DPVsYmxLrC3
pnyBHsOhiVFuEAVNh06yR7W9N/mxnRSI+pNFeguNuQfmI07qYL7cvBHBVgx3QGXk
9p3qnh8j/XByY5U/tMQ5c5B2gwmFWnfDXUYvsZTjIq5D/7WuMHmDbUF80og5fj0u
CciQ6WK1U55yGhyNjYtrB1V230x0pc0f+UHQkpnTcx4JW+35tQv1MFcdUQFkAyIV
ddRxGIFjPRfvayeTg/VqEbErzryRHh/gXx1xKvZKKD9FvfEAM9aUv3FCkn8cNOPr
5yMGlEYOc/nk8oz5usFWzdh+lo1kclm1FxBRY5cwjW2vyZ6fJEDRmOlyW1Emm8ql
KmLvDqoo+wm8IzsdCpOv8k1IHLVZX22qE/kGKfdo+guhqRZFssq46Ty2E9iYWAul
EV5XZwSe39endDUMUKeSqhzQjSrWz/F9yh/YJBUVCeKF+thvVkAGQuqK/xd2omDp
mPhXZr5f+laZwjJ6WBZSj154YaCLclnuu8K2/V/LSw9l+PVmq2zutw4TYwZxAT6Q
5haqmD1ey+5u80VlyLCWIanU3XR1vAYByDfnij1H/rjmCW20V5IZLvq5bTKlQyn8
xVCH595jUeFAJksD+puntK9cBaFdPpOvf5xgKezB9YTTDX1m83WKVKcwFZnttnIe
vNWqCrHBXXQRuwD/HWAbQCP+/sTcEQlrbpwCnDDNAE2HTvruHd3O0GfRQQaPxRtf
EXdHp+59dOMZtPIC7LnaXkBTe04kLjuXIQR+2IocxcPRWqkJdEmLB6F84FQrg+/p
Dsv5w1+PUj88Qg7ssSIoUYpujztECOWauPNRx2nu/OvyI6hSTSI//6SfcojJJm8c
cehkYKCjWQdXBVVwk8u+5Th7P4QwTBoqGmF9T/S4ZFF0myWAQLd/oJpWtDUvyrP/
OEjpdsBXjd2GJoqpDjlrmDUTC2dLxQsCE+/bgfa/bU4XoBN+ksl2JSebL6hlRPpn
cMRgvfqFLf/h3x4P1hJ/unloBNaQHlVdcajE83vRusTOgF3gXEDSTdWTlKxyVk7c
4jej5UCAd1n/PIwmv0ur+OwhU+3aoyrhXpExrG0DKibrZkXVLzRYMEDQMnuUO7A2
kXY2BzTx+MXigSotSaD5Y+BylGYPUY/kFXO0Q1B6Qtu7uVolrIwo9EAK747kGFIJ
eowf0UyKYGh6omHQNdcD9FqGRb//X6ugGbt+R+ENqIvO/68V5+LFDzkfiaXEkpz5
8RGS2EzuMDgfPDI99RuYDFgWfnj3ku1leUlffuC4HB8Jvc27mCs2R/p/Xh68yJIe
QEjeEwEDEVPVvZyTxWv5celPt6SKdrgkETpOVJmmDQqUoROc8bHDTFBQmREAMLyA
T5vL66YYKzHQGhX4quyn6mH4K7m/JArIScXOl3JZ5A6xP1twgj6vCVQ9dXd2GvI7
dpFx0WDE6gHvvvRzDVYWu/826S/RNRMOKOxiM+LjGrmn+t2Q1XSoGcVLZsKcbOec
rG/9S4g9gdqRuE6xDG0vbpD7bNPvCmR4+tItRli0Nzb9HsKlRZA8ZQkzuyuz1qS7
z8a5ZhxF+5Fk1GcWp6FW5z7DNyEa4PT2AM4CcSjNOKYH4YefZClVcYV0eybJehi0
eKukGqrsGwSb4GBnJDF/4eg282wF5rGy1R3AlRmjCG0l1va7KdmcLa+19Zt5Fwnf
wr1RN3alcgk9Z0r1GZssDx+yNPl5mewPz4Liq9ZS5CmoTKumI8NWwa6r/4gTaI54
4LA5a+LKWVA1kMw8De3b3iTzwNAXbLVxHJAvAN0f4yOIdJMf8Sd6BIEkA8IvHQNG
6m4pFgCVaNaQ0c9qgTQUdOK8chqo6jTKxYWMfXWJZA4qyUf2upZ1pFPd7w+on/UF
0DBr0+7IxH3dIByjSWT5V9yM/I3jT+4wmlyspTCH42NrPrSkAy74jMD1RrgMUWao
u6sCbPgGmxpKChJCYIhRNdqWkcyOMZgDp//4sJsZW2cN75nHwF5g9JgBYqHiMCA7
GmUrTdftYal6G5jndh/od5cUAN+Ib/+FcLqIEofLXL6fwTXcFRnIzcNGqkCS2zXQ
eBe8IksCg+X8/yOmUAiEO7fFI9AOYFygozSzsjSp8x2YwlaV9qLU8uz3HWXq0qde
zsDARvYm8pydfPHEE+yvJeHBIiTk7LjqVltKScyVRKIOgV/5HdP5igKbkl8qpLb5
HQgOkvrqOcSsvibr+336Tl1fSjeWcfcfM25DMaKdKIn968lIArxgiEWD96II2qCf
ukBQ5pCmD26ZPW5Hf4KA2ukPG3GXxW8DdtOwDOh86DCcxwZlGQqjWkpQVrSAXA6k
c9ic2bAcUAOa9OwrrgPp+EXLLIdnQhIjRF/lLV22nu5iMzmOCLbWsj4HgNdyNGNA
cWwmgCSGNxOZYBW6kWxbIcUeluDkWlN+p+BK7KvQfPYGliYEWaTkLxVcQmKk5eHL
gC6u6LZFKh5yeaekmuiWBo6SbVfYrmJpNhdukPSeL5SRRi0LqPfi7kiYcpYfBS1T
14MKkQ2Hv+KaywBg1fNbaIaNBI04emRth3CsoQ0uQMWrGp7lNWz4dsj815hhX850
oV6fwqiUc7LGMhALLr8GXPlYmVB3z7yQLEtkzmd52E+i4NUThyBlHaHQPSIVaLg1
ynt4wgG899gpCyDzZQCT25hK9yJ10lA3OGZBwWeMOxwPMIl7CPJ2du6ivpE7dJsB
HeWVukYcgQY3gOIKydc8XFovrj0ZPwY1vRI9yXIilBiqGWu+vkXOAMy/kqBcfK+x
hU0WmNcV8pIXN6lqQrudyudatIP2unNSEY/59XdtuHdS/8ekkuzmlKDtX9qtlj5P
xofuSQHj4LaZpcPJU86n53GrDuovGCIZkXAbKTfx5A2b5Or0ri3g1uS2OXLLWEJQ
iz3+dsLabdJuPCRG+zjTScf+etWDKI7VK5/DDaiuixTenlDLfqZT36La86t7GHfZ
n0NNgZrSMEmatIdqYCGKztgwUC6gQ/MBJA/SO8C4jji9BOz6NaGKykxi82ZcQbqT
gYOsKuPnmMHFh11zNLRglI1adL9GlJakIfw4vCbskwkqOtMHfwVmATPL1XDDlENN
wfIiX0920zjj+oJWjTaMg3v5Z6Ts+5Uf/Ln+STwDQ5vXtfFQgEq+7VRiIoFhtc0Y
6GkiBUkOQerCyOEZVv2OBVWxNiYfh2pn75NoPJ4cG9PMFyAqDxgPDZrktihB4dU7
QTIY3xA/Zwo8OEm92R4DujU8XwpZyAs+4osD5i6FI7Nosb3FK+2BA/2iTwrYagLe
ub2sKFRFISswLO/L7ywNDr7m+4wZdE3dKfe4EfmWsVLqJ6EY0iN7xDz1Zs0NeXy/
xzcmkPUVT1CXR1yTwkSJQCyVIhBBai88WovrdlR0Jt4+/WU0CFy8dl1Py3IDmKqK
CBS4PH5+zzuP/1eBUmshkbfh++ryH+7dWY6hShx++KvxPa8p8E/LbGFke8S7ofLP
Q1KcE0r7IOtiNIt1+o+f92l3wkwctuouxgxTBkM+qXX3H0DiIvnxxrrL3kPGRncm
DBWedEcAqB3DCDUInrEBeLx8BwLf7KqkGhluhvbTHB2JiN4xzf0pUmm8z3BUXcp/
SRiD6bUwpANxdgCDIeMUmFLhznwwxauUtncl4x0fBdtLDxonYJfgGDcB4gkaOLP4
zlMYSgQcQFMnZbLrFb37Xcsci58uM0MiVyZhVVd1eOB9dtqXvR3EIJFv6uOXOca1
NrX/nY6Ve+GYH+2UIMGESU5TbNrNEgGEOCGF1FGvbDLDfMSe1tz4Y6sn0g0R1Zwe
2p7N4VNR1RSjNq9HjFTJVF2FlGGfAbcj4n0aTdcalnffPkyvMCkhO1OSwNMji/0M
32QhLy5sUrwFCs2n3auYoye+xbmOKlMY5uSXFUv+RcnY1Wb+1m7yS7NuCbhn+pGk
oDPcl6WQzVH+9x1Cl51HJsd16WTMP7gpOJNuLOdo8HnnvXpTAOkLFMS18uavX83X
lK65TSpdBnlfDEGVIheLRgMkwsNsi6xfvd71x0zS7kFbOsSXkD3hx2MZzpQhF1oI
324TGDYAs+OMUtmTSgnYcMnvNdahVZ0CF4NHi/VFruskAypDGd/O9udwoGg4UEot
ycMs3guqt6xi1j/jO9dEudAjRHw5SjaAPyXsAvzQX/h+S18SFOwdEDSgdJA6Uebx
tAALSyA820ZZraPax8/kFOx5l/A6+fTEXDRwa3ODrJhvf5yEm1yr9jUhqcV6wWQJ
YkI6HoSiyJ3DK0gh2tKqgAPy53i2ABZ+WIwVlaV1hyI81vb0oRfSWPcMOzytTXDG
zYUG6xVB5nN9IZNsOpT9cuYxqzxZXo9OYIdIoE8sDnK4TaWnSZ3TwEJ4BLd5By3X
rusfFDodOAcRO/r1oxOzy7yhnM65CNkBAHVWAc39bct2DL95Qj/mErpF3u5sfVfp
du13RJ/SqUcbbwQI9mD65sl4IF+9dlNrOMXzAFAz4X7ZhJXOM6H934BDuhMRLGJh
05PMIWkjerhzJeI1TNz0JOnGGr1gkBf3fKNcB9HR7niiUjfQtPioTZfjgbHdtuvS
b+yUQ52x/e/lyRF52zC1XnWl1wWqg95TB+INSKgiTZLb+agP9tn89ASSYDDwsoNe
JsV3SqcldxIXVV40h44oC+84Cul3RL5kmSHw8mMHZ7T4DIMGcKdYlh+L+3OVmTMm
STXa5jJk3KIUvlqKkLmbjbt48LCNDtIcy/aUR+1FQKMv97o1svtpo+CRQJLfnZ7h
a+h33DXo6g5Ekb5MmEFZf2PBmjkaObkIAx1TdXqe1pLkNv73AxH/bX6es4/k28tJ
+CtQErPtQIfN23H1WMFGqgM/oxSshFyZyq7DRXyxCWsNvjeGMqMVra3SaPeDrBqF
h7WVZh/faaq3qhUVH4a4uuBZ7+FysrPDVGmxi1OHZOTmXXpd+BEnEBcVLCj2UZRG
TK9RT8JhQU/8Rna7x7T9hH//v2glNvleDMxD9C1d8qCPqmFs0J2o8rhr+3ReNJhW
hRDzCvyF1Tkc9kC0/PbmxCeuNvvl7UEU5Vvz3L6uJmnxstP00keuN0OSWVgQ5AF1
pwbOW104QnJu++Kb/NJgrggmvQPJvkXfTh7YNtCNKT/1gflVjH8tfW8DXywQRmpr
ulEAKgxt9PzObADBXkiy2gOkw0msHpKv7YHXApX+lv6ZnOMJHVVtmXqfhmrCG89U
4X0Eqbf1cB2F8RRc1/eBQoonzkOlDz4yybScqXOFDuYrgBMp3NXJNWf+79QaAuCP
GEySDIBz3qQ+wwqlnAhmnij/c7aO5g6EP5oyOSLPhtg2eoQYoVqlf35dcyM+SH7l
v/glkn+yl3py/rkyP02vfVtA4FO92L4PTTBJSY0Tv733HCYv2aGJStQcyTrgHt40
S3cEHWpb1ysAZTrEmTWWjkRX2NWyNMhVrxwcef7n8af0Q4L81FISDtTgnKLPiHF/
KLY+JGdM2bSYvCE0S6MVjONxayoFcgfELLaBbvqGFK0a4QUOELDwOESNZ/otG9b6
MrmzGPzWhcUFhgkCux6AQfafmvGLZAvSD258xfQtdtaw6oYPlg0D75CAhqS+URst
UAaxntEK+mNzrejK0+/w8fa3W7wRcpkytqGn+FuzB0ym5kOclLXHYcB4+AR/GcA0
0em7QO5hDYbQkZD268s62IM7kkK43ORtNt2ee2eUFvwrGDkblEeKay49CWLV1ZKw
JG2UFMsO9jN9KDNEqKo0qWIggY1zA2sH+6R8suDgP1W0k1/B2QfTxf14YHmBcdL8
aQAwwL52SC24g0PSYqKwR0pdT2mGFJbswGbcTXj+2Nr/aNOAYv9k4gbq4doyhUfq
H6Y2SBZnWA5MrMIx9i4E5PG1pYvaV2UfXFlKj7wlE8uhHK2F1Ghf/E7xDIJdKP/b
iYK34dTBVXqEEK6lFuUFpiIMbEdQSiKWkUsEkH9vBghU0jbr2Pr26aywnIxoQkXW
imEI6+jtBdnepFqjiixk/k3c+7np1Tv3THZUq2tAlAXe3JEdlpdGEX1M2+yux0ua
K60Axzylvbv31jul6ohMRV1OKG5SdDetRJhsE3hR7k1IKuDq6SpE8FvWkM33vzVN
Bo9g8h8C6kEA8S8H/nNOmsgOrFpdMYhodIY2xrlYnHh0py7CKDxh0+GtKdNbq/KQ
kAvET03csB9VDfAi11jPRMH6Mv1vPWZjqCG9ni7oSEBy5gvwfSO76oGpxO0/25Fc
9HdGYloJtQkseqYNihjdvrxTQu2UJ1MMpZk7McRTNPjl5X0m8NFBxwgtDdvyaAeS
46OnHrLE7CgY63wRWr5WD97DDhySNxt4Jr67UJXjrHx4mtU15J2HNpNUS6gPjOUV
uJea7ejPahdV4YXP2vcF0pkmIQQstVWhxAQwuNLICt/hcDe0A2hx0nY6/PCs5H0G
VjrZ42+lkK9GtiWwxm+bJB3R9Eq3NrJP7GPWFCWryPB0OrGPXLqzwoTap/D5x5CU
SrsYvVqgm5TMH/GOM9FNm1f3VO0VHPSW5k2lNAhuJ1YORIfyk5e6MIBsRkuYQiwR
IpHvuyDOEBO2O0Vu1Wj4PPtHnVWf3b6fO9MmBZcHwbOlygI0HXJwDj4N4AEZokMS
KDD4Thxw+7FzJNACRv2oloLObDOkKWQ0849lwarTziGSkBP6I7pB9iCX9P9T4c6l
FCnUN+1ZsfknlmZKwgBhopXmCSgZmE0MRGlE49KpAMrgARaV+mQOTobKuTVVKvac
g5nwAnG2aU8n4VbckPMghv70qozs05vQeCeLQ5dSWSOEygWKvQDElHIItScfUY6k
ibcK7VFYxWcVQVpDmPKSwKS0uszUl1PW4GDVaqkCxGBJHJUStAwIdZajafhDQNXd
39wgUSbcemnIj2K6PSdE6Bd4AywyzOVwS3k3QOTdCpKybtO+ZeKdHUSKcX1VRJr6
m79otO932efLafm5ACh6iOAZScnraP+cpTRkFfLjfjeUezTRjbExVf55R0lfAryX
+2krM4y3PRGsOjfcLiuD/a8E7mrQ9DVeqo/5gms65/ZghNuD2J+Q+9nDqwGfWxjF
nBpfqLkuAlSEvEjO3qNTLGLhPZ9f7zSKvE28IF6m3YQjIfrx16Z5zoTjFe6iSf98
T9pQ/d8lUbLatL5vHIiBtrxpOU6LNc5TGbJmT8VIuBm2mrz7d8u0A4I5cGhpFskA
cq4yBLAAtAJvJflqAuCZ/O8lrBIhhNsTXkMskV8of8y1ZRKZPunRTCdTGdipVAIC
cI7G7CijEnfkBqzNLnptOK4N9Pl84OZUQE9wcQOTfwMSQnLDno7fwASSNxxOmL4k
S+gogbMQBaBWfeGpLRlhmrz8Xum2EhzSHL4GnZ3cbw5poOzGZiAMOqDASL3FtYzt
I6rmgNUj3RLcabaDmpEPaGBJrcYFByqL+P3LW0ryEdiVjwtcUvnUI/tt6nlqr6B8
x1yPmAEuxtrEPG8wJqe/h6Drp17dKA0CBi+ymal2GZNoq/XHZZ44AMJ8NT6AbNtL
JIiFqDnf3dVl6XUHLMWuJAnbeaJ5Y0VNzV9Lz+qbiRUe7/r3vDDMutIvDXEurO95
fOg0bgdvQH9XLmz/xWrbB56+SReEsk1ZFFqX54q8zX4aMBA6+6g3EjpOsHpsUrCm
Pq9ddnHoXKLeSSTll/Pt4X3fMD3K5lCNvh7aptEG+2Va4AKoQYUNE+xdlsuN14ts
JQwP5Z38SL4otqQbPvCBVY4PllkTPz6+5ZWLspF9rzSmcp4l0LNAW/ymrKby9elu
J5G2wDQQX5/npW/F5Tp422iaRs0ZzudVWr/iLbW88sMv68gDj6tlH/HHrgjziZRo
vwI1YDB18gu9OpwB4r/e8cq1BHzL17U7IwBP4JZEGHw2v+HzgxIu/h10RwAEeMsQ
OqDNd3Q1oeJg6gOTzXnTLsLQ+hlYVKks5cMM/Hw1+vyx8gACufxQ6omRggLrdgp9
fBPH3KkGYtFeZHafpkVvSHqCj23SQJgo0o+hHQwfL1sxZPSab7XMcwQoBC7oJ249
VDGhpp8+r72V8xd+pQfY5JwOo3+TSq2VI/DS78HTcLug34BnL+khXzrn5/NN88Un
DnlV+RGoCpMVjm2iqmgPKAlRoglMIhR5MHhQ8hj7/DUNZKRGGkweV/3P+RAQP5dt
DTyp8iw0v1H1pgHUbQEWaoPHe1s+OFOi2mNDFfA7iyGhYLrEYd7QHmkydj5k6G+z
qsbyIkwplhQPCN++icsmCAHy5CaLTMQuUGZ4iyAnA957+edg5oBXyp3O1pk1vGfl
X81j/NpVI2qh/7JtNpWgE+5F6pwJ550AVQk/VjkCHo2URkBh+630euratTahClOs
CF2XNx6inpiNni541R3ddOaRuz88TLJITBPxDZbBnfIXlnsQ3cYsJPdlxA1iPj0z
ss3nr1XaXJ5rVA4u6uQNW2WuDxhQvIkUVluEb2ospeEfVLoBJZF+pcCjoaZMOWJL
9KGLSVwjGJyhQSpcMDfcNeIvG2NAbuRKs6ElnCCtnyUjRV5VEGd5SZ5g1ZN/vD8g
oXW2vxLvQZksoKrATLAtxcvGQUkqVTUA3iu1lDLFo2f/ayK29Xib2pC5LlGaI0qw
1yZYPwJHru1Z+Zubg7Pxi5lyTyyLsaA1WOQ16xMWwkeoT9j3Hl2F4YjLa5BU6N07
NE2ciAA9Fik8AWsWyvW3BSaw0e6ek7ukwJdfHkUR2aZvrNa9ELrrlRhqGGgV8orX
6t5FyxvkyLRtuMiJ6wtuacXtdsqBHQE1Icp4R0JDgRXyAgl5t5CORka/R2CWYJCw
qbQJ5c/4NhT3IwXs6SPFWBauZcre1fOZLDXFb2mEdrm9j1OU3FVJ+n0tco9PX9lS
Jiwg+GRZiS7y27sZntXm+SejysbnoD+HL4l8mOun81k7cMQ6GEAAz0Fyacg1OxTY
JK0qOx5CzhkglP/pJERUnuhNFI0GWaXt0JDaSlzTkJD16IUaohymS+rpJClrI/Mh
0aggI4EHH3gNlX8oB9VH5Kfkl8p/QZUE5bq4MXw+iSEJS3We03YkAKJg7JUCbR6u
vPE1CzLtqQmLeHoQx8BiPpLhK8f5kj9fMF/6J1xniaG0LpQZpn/g/p64uDpuW5Y7
+RWXOYDszeW1ec6QwnEO7WUdMnFzVBjdVe2MmmiX1LL4CiJ4yqtK0WpSK1V1Wg3W
8ZUJajlbySfApkXbJT1LakhVCCGMg1eR4lGhOwAybEnz+Cs7pWx73SZ4a3VEweOp
/v9wm6FTKlzwyHPSbkQpIZ65OIAeyv+YBOzSVV2NFaMlByCa9b4X10yO7lnDPDiB
S4mFODRRkoTyQMCejqxOD3W1Fl0x4pgRLxcGV6qX1zbCiTQmIh3OcAOMHc82reHW
b1zl0kBT7hNsw/FWQiAaDjX87a+isvop7Y+71VEQquik4bNFVjN1xnngv6mzrf8Y
ji2pIdpyJuVYEFYdhli7E9gP3vldb9hIiQozt/BoBHBX5RdaCZmkTZad5/l8xk1c
uj5dNh5ffsx8s2iyJIy6N5BIOwW8C/pvv9dPy2wHONuqi0KJz+bie49sJL+W8wVy
NHCgXGIGsUCSTPmAZovMU+COM0i62++0mz5b5tcKewTq0ktlh4dc7FqlR9TiPLmy
LQVw/tFcDTTztGVjWW56J34AHZKl0OBIlPzpuDkP81L3FUwJIE/6lWAKx9KqpdVh
8G2JkJF+XeeOLYXWg++sUY5e8f7Oik9WpOYQaRofm0MjMDysdHmdHErZHF6ciwqz
uFJVu8r1yf0lJuJh6dU6eycISEk0Abj1gUuVxNDwlu3xPwna/iMp/7k2uUEvB0sZ
9OjegFl/GAZMdBOOMdCKp96E6g7c1rF4rZDvpbUBc0M0/AJ+dbcor/W48hbRdGF1
iJlHG9AXnz3wFlP+Z6x4BO4wd8yLfmPka1fg0p7lzcTrera1Qj6mvOVz889sMhnY
mleq/brG4js9Wa2b7FB0xUx07rETuhJLtd4YUhiDb+Ymr1VCku2q7j053sTdUPze
jZIASWEQDv94HfUZ/Q4wbZFdBeVQS/A/IE/t5R7OOyB7lkVZkodYLdvAoSs+4iWd
6+qGYNZJ8Qq/JWo+GRKpoReJSBn/oYLMumXdYSG7kVH0pXm4AWX3J6B//AMl0Jeg
NZwuFRvDedoKZfneXBfqyHGXV4IYx1Uqt+TXWAXAMXpZDeH1xpfRyAbR2tGWI7i3
AHqXh5dwFuxegjAbJWp3E0P7COBAUxF/Lrt6yaACWpgKbD5cMErXkuGnAX7Z9CnR
9AOqPUfNJEsJfh0PwTBlag0AEroaNpc0bXK5icN4jR39vUQGLLtqFotbRM1+goX2
e9TSA8OEEA00Zmy4nNxqPWAUeLlKJbLsXogSH9WmHoqPsf1Ld30MRidDjasbK8sF
+8t0W2c/suE/jXBQpWXDjMbv090m6sPIDM289bembCKnjMjhrR5CMsPq2kSFxR4r
AwapSuPsY1t3+c25S/nP3d7+28foZupPdBVtf6OId8NtBAqFmwwkbsevn+F/SEd5
C+GJnS+uSiPXE7FWqzLI1Gz4BjWKgXee8p0MDLuASFTu9IlbtN8b9YlMwoQHJcvM
NaxQnzqUbE5eluuK3/v25dHbSUJQX80xlUQij/jeJP7/9gTvVBTruy1aVNTg3d6Z
IGity0+nl4MkcRKSeUvAVnxkwHlL8LcA4qZhunOJS84cIM4nufnr8LHdUXa7oGBi
1z39F++s6Dg2hnYAPMDNXtQut7QN5TtFpSTbrPzUI6JKv2BehFZK/K9Emw7jaF/B
nYvs4UyTFUW15B6u8Qnv+U71BoyLLMuaJv76aJLmctRLkC1zzyyb1DlU3cJDan+R
gzaoWLs/uhHKYxL07ogA1Mug6ZYz2LoEL1+6BEz6hmMElFcWovXAx5LvIGTaUBGH
OjnNrh1DUmaaz7BCQOnr4oK4RgIP8ccml2FX/EGmaYZ8jSB6KNBCgrYz+X0W54hv
Qg4Uaa7XmqvrKi+dkXFNa/mQGAZ0Jyr+YmKT6HP4HcPrUwMgVA3/n0/tA88rEpDW
9GxgUYLoN45YrXK74zzrX/3CTFIKpMQ25XdmntruPQTaCc44xNj9xy7u9pOXjSwv
JbpjTnZISIys/hau1kBT+MT6Hte2COE8H3QVgOKyeYZ04+ie7/k+luyY6hrRTVus
/Cw/1WUqX34a33FogaAfTVdm5ITqsR8JwdheOGuBEMJZZrH4nVMeo1+SqL/Pz2+r
H7lXuymywgNQGgLH8fTcH2VhyWR88FoWRhxv9c74fD9LLny7TnEhbfIrS7K9wNCO
c27VtJyo3kNHDKYsry9xdOunD2u5214YBJks4qBkdlNTj3Ijj+79qlNDWMfR366c
WSsLBavcFifcj9ZUNbKUoqmC4+ThptOz8woi0hQV1F8SxH4urOvRzEzZDSgf4/4K
ZI/VoCdV5bgO9NasEr0RNjLY5l3CjJkG08TFSV5qVImQ2Ukq9wL6eokCkK27kFzJ
X/LyaUWmu3nVY+nkmFuXcSGk7xHFPGBnMwwQdpkptokOrUh620tms0CNRkSKXvvz
xC00gMzOx4jcIWVc3V2wRqkZ4ov39C4Pzakr7NzlsU3Z/ScLD9Sz/0aX3Yn5axns
mXPR/1ROE35FBJNBqXfP1jKQ0CyCBvw4JcAKGDoMElvm7G3l0nN1HPWmgVf61b/q
klXh6KbkfDXBfrRcNDc01osNCAsG6oAutpjmdgrr7mPSrjzrri3KGyKXyGGYpPIn
2ZTRLHMVTJk2FtDor3RIqIUtnYlec+nRRiu3V9o5xl6IqUB3mW2aIAnRiFhDa4J6
1FjTg6Dkzif9oa3UMPJg03RbHLB/eJvXuDMiig8DIAmDV+QN/yorytCOhwMqzS1G
0vbuuRIW4nCl5tk57zMlkdEdXT+ORSyrTz5Z6G7UrxtlGunZd84plVC7HC1t/5Cu
r7Dcw9pcz0rffcXxGXXbhqXCUTD6gvWKy4shDt++bnYSIl/CdTN0c6UzIwemcxMR
CsByiqJVyXkjJ5+Qir3WqLS2XoBUg5SVcT3Yq5UxVg8SPCF6dKFxxUufezqi7eRR
0RY0OHU5DD3CUk+OQ+z5ltFCD6nja8jUilsA3peFLt922SHWs/zDf7tQPYI3ki4L
+6fEvq6gsKpke3aBdZb7Rov2bJTomKvB554FoInSee9na9VDUs9PDZ42QuKU04wF
amxKGJsHAfJFw0HQFOfLtkQW0CwnQecDdFv90U3ts7Qmsan5o0rtAAnICnMVSaEB
Eta058h9Qmc1rnr1mtZZ79E5V3KIwVlTOu12ikDt4o8pn9UMHAM8W5PFx6NEBe6w
9kabmdiZx8mXSIgLC2nYC4i6eTRVjXNX7YdLvKW46aQAKV7zqIi+nKkrxRmXZK9w
vDfxfpGpP2J/abDiHBDWtYBVvPkea3J4gWYNX+PpnqoGMTyZzd1pEUwD3DRtHw1q
uLFoJbu7Lf3k8rV6yotkKn8ZNKCKZ34kfGCRb6biu1IcpNE/J5c3rGx0HCGGvk4G
eJ+j/hOlk2zGqR+fRjgSP5DygppFXy6Vqezyrc2Yt/Og9TouSBeZpfKqUMWX8CoE
kwQpcMXhvHYz8mkMkMAc6P5ggpNFFN5sOEHdKEFxxryFFahNRNLcaVU7qqV9h9ip
ESUXgAeJthuV5nwKZhxgDdn5/FtpPcHFwA/n+3RYiuwqOymMYRoUlytXEKJjTYDe
RJfTYgBx0mJHzYozL9FC4q7J5sBqQswQLMNQFCphe19lCfi7B9dbX423p71/l4g0
oN4B5CIVTnqSUojJdueuZ4/C4UCAfEGBZCUHIHNPBYMqaReXz0shnKTP0FK92vV9
vsb0/IdbVKpPSRHUV2if7EBPEOsU4QjRrwktx2wbt4oUACapZo1wMiIxpTlY0Y22
9aCvygbFnVcpxEmUUXW3i7cU6JmeoTqjZndcPW8GFBb8Y3VxzHYSVPuCXlf/5ZGU
ne+eLQiK3JU3RHkaE3Xd/z1cB/zJD6e3qPDgNZckJbW1XTO1WWYLh6MSgBAKpgeK
uge1DYi8cIf7wQ3Mk01gM8pIHbFv7HEC1SIUVZfIZBKlFxQSNWjDsLqMuU1AI6Yo
WbKtiS/eU85x1S6qYlYQeFP0s652jeRKX+1vEXV/A8enCxa1y5EDqn/PTx5FQWsS
YbtsopdvoxZ/8sdt8QRCcwKaMozC7JPrFk+Y30FHrecTHhy6ujeO5KkE0mssQRg8
8FKSVDgUdHdD/VMKTgucSAYfscoB/i3MNn2kDCbnATM3smEXRpGdNCAwkEoOyZbU
Js2UeG5UCMeg1nzMzcu1LlI0eotVJDpFDT8jZffomFi0rKFuo100Iw0Yyn90gtYE
Qsn7Af767d3yAOIWIqso3Re2NTIl7gKgvl/T+2YPYjFxDPKpEhE+2lMuB8d04Fx5
A0AoDhAyrwzvwSMGRnBZ3t61XpnJBIfdkOUz/n9FhgBMqo4FECT97SMhfgcwSB0w
oIxA5EtS7IZQECJ0fspMUARJY3qYX6+FN0yMOZjV+oGs/t/0b/dHUY//8H8tbfSp
enG/hPdL7tA4RKukCMxxph1VF3w6bgYTXydlgYvspHXpOnP64cY9xxVCOA7rfYBO
VA18+AJDRiDZB79ZuD6lCgdoh8MkY2uul7vJVJ0NRkZTnOviBsfBNH6brKceNGLG
2/vktmwOYnPPt5gLgL3FDJGq551WocLJo+rPxrP7x64HUuBhA7tG1xijOmGsf45Y
RPnJ2/TU88wcW4wk9UVFfZ+m++ahyn7WtJt1QhtwpJwf888CCcMK5hEilaz36uE2
EfCo+N8iUcUywtRPh8Ma8wlwshPennWckhC5SK7Klrhp/WMop8WbzJboRQBfFM2m
YjdexbKrevV6lMsT8ClHgjI3K7CV8eoE1aAEBXCNWfqdO80yPgnCmN7waQmRUTkf
VIPrlyt7XAGIXUqnJnhHAyfZavTi2KStXnHE4fKiipxGx7cBp9wi1qJuxSQlz+HF
a6lxEI11MYnY6jcC9cAlHW4qD6UxZH3/wmW3nYvurJgV2vENolH4eGvJoj1dfo7A
pLGPjH+K3+29B5jqRpYHGvYTH0NxIT8NeQvYqptq/D1pz5tS9QEOFFDJfwH+/Zjf
HNfAgO+sWgjTV9Ri15t0r16S9DuXGUma0k8BTgtvSeekFPtjKnY+I0eM66BOt5Ng
iMNFATCSMg+gKvlTsGE/BXcMGdpPJUawMzMQJKZYo/376YLlmsYj4mB9YX+lqQPQ
D/pCA1FJ4OZ06jefc7awXjuNEPRHc/tcMB0kqYl7q5DkI72JBi5TeLf2m2vdtFyh
w4XFGwK01d20t02KoySu8VHDl7QVuyp7mecXDWqjvzHDSXAD6OqPwsy8Ufp3q10R
U8ogtukIbc5XA0ew/LUjrovZnzxp2Ds8eIWscDO5JRU/TyDLxwXGH0lQiGlQO8Ij
m9zyJAHVmbp3WxlFpIIXwZNbxg3sCi+bCmXlZJsYrHMaoMQqyBQ7LfoPcDDCK8rg
iwfwPL+39K8bAv/ISu1WA5f04xLMYJV/bxisa37yQyqtNAACKQMU+w0KYw4tThS+
3++0NQSsB1ODqmtbHBlz8KjlHJUX8IkMt5dLrv7b/xLqrtMmGEH7fGtnXcFDBlTf
iyy8AwIKuvrKGJKKw6pfPBaDIjC0nsnCGAJ/zzPzlBCa1efWWEcFb+KEsT9B7nG8
1BnA3ij6VUwBF+ytR+FdcffitHoauiIrpaLMGjyUI6sMYzKuepH8vPR/fOv2WQkw
+ut5bE0UGmpVGx86AwzJ7ps0aP5bCcM0M6dBuJdfJvEo3VQ8ApCaLJydSs2gM7cv
65zMfumnk/6QPmNfkXJ+3saHMqkZX9qgu3mbSe1/2D4yVDKg1jM+QYKHKl2tYV3N
uX6tIE9v6X4MpGRJmi23aq/GS2WUNhpct95pB8SIMZtvraNFeIrR3tlidCUPhjEY
J3KNEmjXaYW5L/2scQMuG4DMO/ntL5xy6yNj3LL2uzgRuMAUClD1QAR12eI/mNZA
saTFYo4LEz/YFQR4dGWUgU9I2YeEAOBBCKV5fBaQPGjMMQ+4WVwnzTOPjCiK4caC
GEtdwve0XZTE18bSNfIrqGH88qj2ULsL05msjTd5jJ1JGTCyO2VCB7kGXXaUI7zp
CMbujN9bUPJu/FjCJM7FlXbOGVkXOcVshJ8c2HP3putwyJWgD6w+st/Z6+NRv/uJ
1PDS2zHvvQlDhunYg5hT90WAKbANzntTf9SORt9Pi2sCDLakpL9nSandwuzrBaFe
a4Uc+mZygbIvrT7XcfTWhN6RGZktVNELbBd8BXgwO8yjhr6pUQWx9lHAj1EgzZRx
OU5A2+d2le2yhK4HqUg+8PLt+1jG9ePDlDXSbUHXiRzfc8wvr4rGlCJGyNjtVLOb
oL/e/c6e/pWwFWzIrUaAUFi/mt8GBaDseWqeYlEOybDEUD1ZT9HLOudCB+4tquFg
SXZ9b+aBzMxLdNLsWytZFhC23t/b9F9OGhLQ/yURkAUGLVLMFTcq1pAQK7Sf0utR
ciDNiTLyyCdyX4A2FunV3yEokcd1Yu6SNRSF9dmI0KlroPT8YTwcbDBpWyPaiPWK
5qa8JLEA0iT1ffM+9cEXJbp2nH4iXZ1Ma1LWUeSj9sOlkua8h+1dve7xtiNQFAn1
rmfgE4k57AfhH6zoWi8eAcTF+PTuF3vq14TA5dUdgCQuvT35TKYjazK+mXNZq4rq
gs6M4DuHyHsnXh/1E5RwCKgWpb4MXbaCe9w5M3q85FwKf1NlKvbev6+n8EE0Rzbo
q+N01mSmDVBKCJgUuXY+7kXTUu1VuaI8FOtV1PmzgEwSCtfWIV1n+NzLfRcae+rf
tFwBo7vYwT2Muy7qeIdUhAraSFuIPhPMRFvwkUm6GQEGHxHOTSd7jK6tRt5daXSd
1nfGSRnpfz3OE1zr+FA0RQwcZ15Ze5gZRBmgRB9dAkY3ZlKPAeIzeHb0Q8rAYP8+
V7Ff9yacnD9lKnLoS2rHQqiSPQyvBanfACyUhhYBa9iOAmoFLJD19goD6oaXctZ0
uwZfnfZnQ+FY1B8QFZZt4tWadnlXD4vrvQWlb28w9093avGLRUyyDY9VvXZiwJrb
3dAKE/dlnN+cEUfmSabiUT6ppexxgzSRmPESvrLRSo0LmhlwUlomgWGCkkgkFPQI
OmDCjKaHg1xOwIsUue78Usg+NB3V2UdtKbp1ivtBPdsDIBbm2hxu1Edhzm4jlDl+
fMONyxvzO3NIzNb5USf3TyJSNzCtOEIlxJQsweDA8OZriyi+Gw5hIA/pBkPyvfoB
v69LY19NIDgktEp42dyZ6pXn7RTq8izpIt/oMQSe5mgejm6dUfCcdjasx/xRzdIn
zu2CRdUADsvPEu4Rb6VK84Aez1hJ2aGxQYWAJM/UuCn0mDnEhdKC2hc0iCLvujoP
Zq4ydu0xn8Mr9XEGlnL/L62aPhfb6v9qdYgUjAS1YPm64A7zAMMnIBZ8v5YcFYyx
3Ua+SKAMNGcLdMmATq8RhFXWdiI0uqXodGyMr4FFOp454CfGNTBhe6IvuZmjCtGj
E+Ep2k5XYhrePamxtuEIQBtY/83owAUlucN8bVEIozlLZeLhw06TInwNGUhgglJq
MJvEdltnfw+LVc7mg8ipC7XuD9GkCGBrpyaPd0eGS1uGHP3APMDEh+x++EKl7Tpg
1L/9vHyO3mHYJET37TnQRV0w3M6P+Il0a74Ez4KJBOAS/ND2iWARQxEBpq1YwvX7
+QlX4d6DD/eeQtlOiezq2gDjHa/rejAQcANcpNY4E5VsWqcOK6u6+AseOoJ7sSjd
KFpM5LucM8MbaxNPogB6EzPRpMysNkk0XViQZL5HVtgKdC6EeBicsyWZ923j/2tL
4tQNjWIKrK/EnVq6wMbBroeXI8DJeOJJ+RVUzpFrGO/sNxvFS9wQXcPQxpaGvZem
2Rux0ODY6um+N3peqwu/D0hP9rVDNrTvDAbWfJcPsVE2HcGOMHd05YZnwubIofX1
t8pJVSJd8L9jGzvBy6WgiyFWeaJM3hHn8yYIS+6zjAYcYDqy2dUmVkfOV79ubf8L
XKHGJmem43NCSGU4bYSTKsbKkBtczzCLuj2/VcXNJ6na17EOCWl0MhJdtTmoBM51
X5PWm4O/1sArjp4x32TMkd7oUTwVxkNN18PPZ4CTLRGhv/UAhfvSUC9xc+9BpsYR
vL/eO6pWqYB0e24eNiIYSycgjtcm5JCnVDnqQ0gEw7maPUKsaWYCCN3GFkqZYmsh
6qhqdfz+kljSF7b+TP31kI2biT6rx+nTr6Q+XnjzIw4pbf44d02PqgGzlkk0UGtV
NYwt7f/RXtA4EjOIo6Kbtnr09+ZN191DHCkHq24Iak3iQeai9VMK76g89Og51ZYI
SUhoP+18DARNfXpPjBCblfNw2UWst2GkI8qFSpe08gx29K0FbRD8joHQ8VGbgLjs
uN1BoQt0bAaFwLOwlregAbdNpme+oQi2N5kg56aAZN3gxykrfzdzAysdZrKgoYe3
rT5VfR4BqqebvTOrUGuzs6imQTy0c/Wa0d1yHFYGviOTGgoszwMK/vPH2yAAzT5w
OGNq5MQe3N/n71xh044PdE9dWiy/ZGGxNveLibNgWyua7rtznrQ3twhAzvZiVzMP
Dy4pIikt+kE8FWpXmMOGbncrhg41CxUpEfIV1+TyuXnDTnBKuZd/Tm12MYgsLI60
t48xeXa0/Y4XoXftxuHxZ5zN8g0h3DSlfsb1hEMeI8AXGPSpOPyxYXyz7sQw26zH
yU1JOV8iO0hpfPk25ZXeGU0CS7hnMiOE9eR1t8Mx5N63xdN8cooB1Zyxa6xux44W
s4yAVCs8e+T4jNMvSzC5tASHp8BkdIncYa07f+OS0J4l3/vaI2hGETDuSwGNTXnj
ah7LSrfyrM+NwpM6JuhjPJHJlifprbLlXm5bYg8LMxPp1tRTw7SDWyoFz2ZmYc4+
LLzCXEKg2iUmYBBcxm04IaMsyJAq0NEVQ2ncP8XuTIUXIhmHs0R081nOY7mt0fG2
ArECQbDnCf6jMnzo+X9SPlfGcFUbEZ6oONGQPqZr5N59J8RAAABr0lGYAc/KyzQE
2J1aBjRgfIJbUuEm63hd8E7Un07rSdrrrfKSpsv5k3dB8w+a0J7Xi4lgQZzYxxEw
5JU2uxDxUj3CC15OhjFiL/Qd6leVB5WjxBLW9F3ZhqyiUxcP0R1mi//jPfkOe6Xm
0WWdlneX3Cw/8R2drY0nS2FOaGSrMkEIWhrjkLW2vDa5kiIui5HzqeSw2zH1VEyu
P1I8eXBZPVjerVL3avi3NQmalBIK/9LNamFIGXsjVwVVczTaOIpKZMIKK+G9kcKF
YxFIwGNKREiv4Asia9ni31Us/tbD5EJBQMvYLURloYlsV0iibbvwYBoyWVeotKaY
uUgnoK74o5mipjfkoPhxwLyOHDkMUyLLMtyG7AOP6nA+pP7ZPcSxLPtHf51TNirf
8XK8kvdLa7YuprGfFd3cV5i5qE473JTIp3ikUZ5L2vbztLfh8Cfa0cGdDPlv2mKS
OFXbaGpBzM64No1uheuiC3a2yzyVEtm/g6tr/KLBNAzkYsDhkbtvwUHtH4ALH1Au
sFz/nm9zExVcKbVQz85M++DNwtSOd+AeXooT35kwCqkeAUEXRDTsAIv3FLvUnaAn
giED6t5Fi01BFSMdSyFoz6TBhuzSxpyzKgr+U2S6W0tgq80aJMg2X/zXBNQebeeZ
aJsRE13NMNbH5+pKbQH4cU3y+KW6JbRzSuFUXTTQ/iK+4JYkya0sjHecmnT5t+bF
tqL9O6vyik/GuzVwrOZtUO1l80u6FqbyFTU7KrpKG5DAKv/OSdfq3sZih+GxGnKj
Zfg1ztF5xoAvMxSdvBNj34nHZHtITPfNqhhcDwMVif8AOtiVHZMiOWL5omyijLOL
PJXn/+tAEq7HBk1YPLhAFdIoD1BpsVBlKYzLvHIzLg4hQOunzaXmV0V46neIq4ag
OrWpRk6CLo33lP5kQpjwNMYLE0J0dKaTYqGqUA3xHCMNa8Dtl70W0CearIVQXwKC
gaLYV5/uQlN2y2dRH9BZqoPCFlc8BsirnAwr7oUMB2HkfQ8QhGOI0s8vM2XVqs1Z
NiQUendIMt4mSEJgZ1BR3z3yW7IIlIVJa64mkjE+MzfXzU5HFCkMJOxyt7+BePcK
a0j2MNYmNw3q0wdQfG4BJj8dRIJFeJgMIYNB9I80/O8xRPhyNr7vilY5shpvwqzt
aoGDuBP8G+YebcWx8a74zfl3MfgXtBgxchNZcGBooGvKFeWH1sMHtXh+S2q2PRDj
/AJFLrLXBF2xdgg+ggEZjGJeH+M4NLFaoyYSka7tBZHyyXyASAGIMvQQDamtwBzm
B7CkjnLYUaqH3gDjSeRyoBKr6I9N+SWIAfiqO8dz6k8TeUamYhsnsI0VGs2nOtYZ
gxLP5bIP6nTaRl30DuMMevZpWyXijW4gU/NTAfvs3uqBh6Z94IdhaOwONejGEpfO
L9NkQU1LNIJMZ667TSiRGy7U6XwcjyeaFgj0Irs7jfsx795ZWZx9kj444L5FFUmi
A7mx/a8uHoaNh5k94xTaTxtwwDtVeYP9yNRwJL2WiEPcFH1Wz++ITWev1mgK+sbG
ZsF2fqaQszxjX/d8e6Z42JOceSrhU3ZKHtgJ5vTKdeWnjBn+2XBWvQ2/Pr6KkKLP
R3YFKxyVAGwBfoEUm7sEZbd944YMLwqXbERb6LJYWI5r6mquRfXqQdaJTg6mMkOl
z2t0sdNQV+DrwN2MCKjl/T9WFUcPwztRgORO1zucHwBDU7YMNBi7x4khXxLDcgob
4MCmPv2C4Vp7J7d/BqdXyMV/IQ1xGorhKWpIl7d4/4CV+2Scb8y6BLHY82PTh3AU
069Smo8ZjbsLxY3LRvbYCqiFfJOHKC69iaEtUMXUFRoLBcCVZd6pbtmZNd0bitTT
Rrks9urVcrBq8xLMSKpRR9akgZ2gzZ+ivjXEMhPhduapgaYTqBoaViG7m4cnVbFe
+9UFOcrEd63kEkYhqZjXSgeWBjzk0eJRW2/FDd3KmLGcHo1jLxTCdNNps2MixbV+
SJPHYxSqos/xS43gmdgRK3j4SvPLYTTXiEdH0qryHV2r79CQHt/OOn9SwhGZYaKr
TeeFN6P4NhTrJU4euYr+479P8xJXU3nDGmzmz4r6EWuZOSW7tN+5dW0dFpr5HwBG
vil/OV3x095shcoev/3UwZbkql4W2Lvyu1pH8ReZfnv9FlqSfkX9LciFwRgndrXt
M6EQP1FFbvGc521IN1x2mOH/aPGkj0xwktlyndx4yPqCBsVHCgD8wqmO52YyRBo3
h8lTb71MSINTEBYO/VeSKWaVE53trJh/AHriH0jILHyGjZQGg08HWBVoDkzkor1G
x/vQX3LUD0PcxrYCXKCBz3msAUK4qrZT+OmvGQO1FBlbtcWLV8lUV54nad8Dc7rC
SX1VCeP0QHgMhq18MGusdpWg5U4lixjcgVRB81R1rqfUJjEzjDFNgNP0H277bxAy
wQUyc5ZGZcSxy2jgHYOxV/dzRMVogtwfZ/GKeUjUPtyAs8DkymLjVhBUi3FCu2II
3WdmTn0dQQ/2KDoTufLQWKH8nCoYIcwhOQc2O0wiuQZWM0lsNLP7kVHuA+ktVWXW
mNMenCeTn38GVNCuiPWp/ProQGEghKjNieS5uDjKS5MmQZOPuCRCeSNcKNlAFLic
eU0VFtsh4RfBvrpG3YBQ3+9OJev6hgsu4heh7eMIvbPXERKdyUwj3i6qTItqUN8U
Fc28bm3QZ8OSFg/98KPK08aw6AdaGkNX1YPNHlnzdS8UQcVC30OsrNu/UfKHM2ZH
WG+rkI2JAIdBEwdLEgE0W3GxlKPyn/God1aAXFLvf7hIX1Nn5wM5JpeuaSZ0/YZ9
Prv/tA8x7DJYg1OwnCVrW88Bxcmnd9rkbSbHYPu0c9zPqsXfBAqRwKDQG/Jx6jyY
RYj/BEC5vXpdrVZhnVtJRUacxREsPLfKMgP6xegiwf3KLqaG8m/xXRDi6G8ToMHc
K6bE7IJqy686+B2IDz/suEO3++dAPoBOP4rU8jdKtcL7/+YYiJyTJl7GZsvsCRIO
HYHXpMTQPAUxJtS6wjnmTdeGOkHGiscLiOu6STRHo3pH6I90N/j1iEXfeZUJE8y5
j/lmWOnq1+MSZU/pSNR9ut4UXOUcyLdYDyGbvYueYpVMCHq3+H98P82mAjCwExrE
3/Xk6eyijdjhWbzyzV9gfJzU/gOybEZIJlL+hXxCwBgoi8OvyT1BzBqNnbEuytTH
H+C8EAN9AP/o9Yls0ABhswEJyTHC769xrQylUQYOP6EFPPPKIKH/NJwi2de5p7l0
xGXrSGa0SM/tt5OTfEJJXVn57rOFS1r30TKjCY3hIQ+gm2Ov7Oenv6fmMvJKRzJ8
0Uf71rtNiGhDgFIk3SixDi1i2U4r7zaCpQmIfHQBDajFAejTCYVR1PqNXp4C6hVX
NXPMeD3aazgPUKAnoW/x7/CVsJDFp/QhCXPH74DeG5B57hZq8Jrf+4R+xXz++KDe
EVp68N/YSaEIr/+LHzZZov1aSCvFNQQvA6n3AkeLexZRBT5ndmvC66v2DncMlz0y
Ssb7Hz2ikwTBF4L6HM/jpQpNWGcuie74BIxWKLnQuKlQIetDR2wWnqa2LjWyvZ2M
4Mv5iFfdIiiaJ7+J4DPlYIZEz4RX7zZTdK+f0nY/TOQPEju6SRlszlikXgQi5oTP
hDofxRBS3eZG74i+DFd8AHomZzc14KsZqVnSOBYw2f7P71KOkpEmIVXOXAhtSpA9
3u6xjqI6QUVqabGmD0Og9noXSuFO9UpahzOk+xIfflsgEe3NtdTKZgy4kI2R0tHq
l5kGeRMVxRoy7cLzdn40NANtlHjH2E3tNE9VoMDJclLJ+tEuI+vrRHPDULw/QoJ5
4cyjmo6rYqB8O+BPk5uHjiwKgkxK7iCUMYO4Te/vcvV/PIQo2spcFlPFNbioNqlS
mTsr5dlknBDBAAtuPHC1ehRyIyAlhy0JYryFLgZH5tdXzXnrIgS0dXvz1UH2r96U
Uu019Cuec+JPPSekHJGybivScd87MVuMDq26aCrVg6Xvl45tj1+OjvN3QWP3fdeQ
OE3MnhS40h3ldbJhzmrCgB7jG5z4LeYHsCpC+HFHCyzSXDWK+ipvJ8OKXS285Ou6
o96bpJ463c7lYhKczwkQ59Bb2KUB0X3WfHFmojtswBRYnEAZXjF56I7uyLZIWRww
dbKxIcDI53Nz5Fl+LWQcz0QbFgPVylAAKrfgmTo3BKXLXwqMzslHXzOG0oZaIqjW
tOphf3WrBADW3+CrrLuHGcv42JMLTPIk6JaDvxPQjaTxd5SLW8jhje0kFzDUkCZb
tSOCwoAe1th8a6F2pGY7SFGFpeUfjcSBX26Ss08UMQq9EuPIlH1KMA17d7tl4Cr9
yE77v1dknz9YeXpkJHSfRSYytwl9ThjCL3VC1TauIZgy2StarBsB3FVu29h8JMYQ
cApNrnjEc8b64nQyIEl6BVS00dkx6zv0WsVzKY7bPt/PhXRMxr0b+BYu8QW0hSok
89aNT/g/NBhjHcvn9L0MDAngIvb6VkDN9v0Opli9ncdnTJpNi4g3lpwFOBgMmhf8
RehCBioyAT9eIvkqK5fG/T8PjC/mlFj1TuyghrVZ2XRnb0+u/JafJCSvOC4oYNJY
xGMepkM2Y/0QbHeWe5Aj8brm1ye+f2zswCaMnw/UhIbz2fiiEYb73BsNa43u82kl
6iyBcIOqSPWKwxWjvSY6VoS1N+zKs8FwjM5SqCb0m23F6tiqoMTUm/NGps3Y30Cp
2CeIm8UTgi6rdUAX9AuO5/kvg9/Kq3B0r1mSuWEq6Sp5NGtfQ0Lg3av+4Khnzldw
LeOKEx4kee05MIBiT0GmIsuoiCOapsKy9r/ILyI9K7Vp82KMJ+virALXYpmpdEVJ
NztXl2n1dYzB25wgpujE1HMgEP18RmAz+GnFfPcpEpogzE+bObemuromSOqCagoQ
O+04eFd9FUDlpS12r4s1bB55iOdGIAdJB9vq7hqY9TS0/Qs+uw6QMiLg/OUxTstE
PI9CHSLtojkbyl3Ronh3AoEJzB7TmihwJNNjD4ccOfEjMMOoMpaefX3AO2vxrWnk
sy0UeiOouO/1sDqHkx8jv+dNDhQbweGOwstt2sq05S7TPiYVH48oMr77ZXSZR5nt
zYlIK8xHEItJ6ZWV57XIHBq28ROePH2tQK48mbsIyFC42oe6E7IQ6k3xImEpSxA9
mk/dr68EG7T8jm3i/ci1/ChmT9KfxRDedK22RHxOAeBdXeboBvA0kEUOMNXOzQMV
5lGSgqs+ZcQZSHsIzP9QEJ+RuKE1COVGeL71frIBJyCt/GlIAVNTCELsffAUW4p+
Xkw34WnuBLCuyYZt1FV0GVVMkjipYHf9naArKlNds4PUAnP4gbPpzjsR+3OPyTze
4otKQaLigmEkyvLmolU6iNTC/i4IT2uxqMsPImjpe/e5Iy2S+Uw0UXFGW9NLTMIZ
mB64ATSEt9JS6VSaGvsAYwLfwWjPp+9GOYiH6Z/EGdWON8trZj9kTd59ZIZ93kTF
Vh+O49HmSH96LuQos9QgB1sbkJ8VxcJXeu7dqAe6x/39WyV66GO0/5MzEQQiLMXP
JvvVbsY7hoqbQCl0spi8TH00+KNsj5T421ZA5/SiV778pmsdW+y6eIQ/d7y5tf4+
Y4VsLVhE9OPiTxBhWges3DQFxKBMXNS+89K+PUT89AXi5i6LtBm+gudCYLAE875M
U1/oJCJIORz4rFIbKOPnSZHXTTABzT+tIe2HmtEM6R5ZIaLocjRFaNLnVCRYY+0K
28orQhcevwdsVt6HKIxA2JsZBniCiil9K0aoee8+SXY6oaMP1d18ZVFOV11SDQxB
ghwwFjwe8d7WzST+ry6iezu8ZXjuDt7YcMGnHRu5DGIDTWIDq69Z9Wupj1Hr4sQq
GyK757WJLUBtrOiiYXSkcMahODQYxki61UjnpEV25jOIkY0uzK4ETSSF2vYKmXfQ
vozITOo9AjKenqygBf9CXOsDMgzp+o7JqYPOCIey+S6oOoPGaZD42rTqt3O0PGaV
Cjah8qqIx+Mz4ahuTQ9XW3OMuC3bABqkLJIJm/LzhCUL3DbrH52PukvKv7TPOqPb
XBIn/7hLE9aCObextieQgI6+4Cqhpo/Ed4fX4+ZYi4IPB94xkfh8Q++0MLCCd8Fx
PefPe0Oer5qts/AvhXHAjPdW/32jbCbvUjKiVAteqLU/9eJRIgimaCUQQe8qopaL
M25Odjl61au0p7UkH1IcvmvbQraMCHHfDi+68eUTNUfZcAymwYAHbK4BHKLn7J5K
hseVv8JxSIiX8KOLl1VXF3G2EspYzAF2PpdO8LaOooPvld9wlixoftnMIVNppnq3
bQcAtg4c8uyz9k3MJMtup34odfZ2MTcgde+4h2MF2wkD3jBfQ3wO2vOOnxd0KNsj
1ngRFr5+30mPykgTBd7e5s4iynK8/35w6/bgHjnpclNP1gHpFdod8W5//9fAMvC8
TAcx+88mKblN5MBvUFOcJ1+tY03D/SX9PF6AgyEf5suFzbYNaPqYwMEHAs8jtOl0
vr7QwSYFXcdYaycI+13b1lDjWTu4y8HxdwrnrC+Npk8/PvpYrbHm+XxF+c4wUA15
Xnxt/x6XmgD6se9s9ydVdUQZsaQ/47tpxrCQwtmRIVuhL+E3KKBWVICA10s3M/zG
/yEkKDQ4sB6Xkibo420oaBN82a8uzbCRAcBDENsP6G5OlK2t7EgxMsliA9ldHGs6
YumCmG5dIOKVcvwzkSSczpwkD8IxOxuEsFiOFRV4ntYV0WknBpSjmwRdzfAVa14f
N4RapVw34dJ0pbiRKTOEAz3ypraIn59JRQ/90VAQLJIF7v8O/k0ll0v4WdZvbS0N
YaGx8pjl1Wq4/WDK3gVXR1Y9Z7LCvx3RHcycMFejLyt0ubmHNuUiDdJzcUZ6gscn
OV1H7dotMdGfv2UMXvwNM0U0+J0WK6eliPpzyMGpvSBDoyEhGuIUj2sJhW7UZqDa
mPJMNHa3ehO+KIOmYf4n4OYI44mJCn1pYfG38O7TrGBUq7OR4bnLDY+YZ1qOrrr0
OdgCK3px1w1Qk+TzdiYqckgo1qPni55xSajirTUYcDPZVi7BFnJ83DWIyKKK9+vj
jeqtvmCpWSgIhlohSZ+oOkcZtNxCr+BQthJ4JII7f2QQu0bNNULavzEGV9YL5qg7
azGftyxru5Y52Y9FWmtIezZBYY/xNhdxbDIdMOIUvfYsanMZQQwVGs4KWirklxA/
pKNUe0l3WJh2l5XocWNJc9VGQyd2YH4SyWHpyUBGOxITLUBqhnBvcl5dcTI2Ix1I
TWmrmy4MX93VYxFTBxgm0ekAFs0o0YD+PDYYpWWRAHTAAQyqrCo3t2Nd/cqRKsnq
WWW5uYvjR2QoBVZpOIi1cDPaD5A5LL50hlbPo/q/Ks3rGoKMglVwb5aM4usDh4TU
tXykZVxiYLBeo3n6+OGsjCHcoIaLIKIg5t+Mbg/n9kDCf2O77DMwzRDstSBUos1G
0x8RoOxxcbvLz7sd+ihlTus/lT1S12TWKeminp/Emo+BKscePp0hYwbNCPdgtGqI
NsUtnzQKPDhJgN9zBT5n/w5Quz951J1FXRmJbqUC4SpBWizWD6FLb3zwPVOQLV8O
YPLyBcn3HeYf4lEGSBtRyGZoBy9NJ+fELv5CZy3qbg2OSnLQLpU+qglvUc72BDy1
aYGIf42PX52IvCbEoAEhb5ms6fbRxZ1yI+13waURMR2NCPC2KRFp3CbAogkaoPbk
ayhY1hYMNS4ofRjoRJdaBxjt19ARR5p7P7nWfkH7M5APBrCCwXOhuIyibOHn5ksL
WWBxR7SK5IwuJ+qWHxvc18I7vkg+1ReEH4DpOpTP0tpf2Bbd0w68kedr23z+T3RO
+XAWdcYeGQBjGMo3l2k18JwgmShNLWkTreVAOENpSInjDMJcnBtl66Y0sh1a/71o
CWupreQnluFbr89L8t3hjgsc6Ea96IA4s6S/I7w6Cp4cQWckla4j0H+v1CxaSajQ
KBtdICs1Hd4gq8id4t03ohoNPNnDp+P8byD+59NQYI/2BIRox0Ug9gRo4G/nwFeL
pZzoe6CtMsGLR+eOf9urA/r19mmZcnh394fB3LSEiaRZw2pmhgwophAIAfx2SL7g
oUZd2UHnwEG4cuVWKA7ky43OWOuZBt8nTKOG2p/pQVrFqDyLfmrMEQrtwIkuARvy
4ves8X7CV1HpB507Fh/CMagDMcqeDRbt/EyvATNd5LLZ6xAzHkZqQSgdLJjBpV/w
z35Y9NbWl5dLxq2wfHBAPkiN5yI5LWxtnIcReFXOG2EMMYtRGN1+FFSz96PGhIL7
ip38NUFnXJk0HecvrekB5HxCM9h0C9/n7XJhd61RjdcYsgeTROGElfEA5fUoKHXN
8h9OALibmJ5UDR49URWt0uPVvlB6UNT7zEUowIEtBsxo0dVfhl0DTjR1OvDvkFW1
uPIo3sTGAXX2YeCQ6ByNKNMP+KYyvL/oM44cqQGLF3FErqRSbkqmtGeLL68H8XJf
SYB8kgGuc4u+uOw7pnRtlStCq7x/Yxs2ZxkPD+ccdIcMLqqOqRZN6RKvi93oOqqp
Gm7g5bjeNY6JmU5AEliIVFE/hqtus0M+/BOtHJuh3lduK9oMWdKApfwbCGLbnL1u
qgvqQQ4lTYu+D7cauTvoMiYoEplQFlN/cIz7N6MvX3Pz6QYrU375v7gCjVt8bbPD
0PuFt93OBYuJP+iOAi07+Imtgsep9NBjjTk2/w584wvgkroNvW5MKyA776Ivy9r2
kNQ+L9G+xwXgaGdT+aqveFmlzCbA0GkuWmwFjMUoUY8wwbmG3G9YtYcYHO+xSiFw
rCzS5qH71WNcskWvJAU27pti4T5uE0Gisq1RfrTvephk1boISNdEmJWqfh4fx86e
vsxHZuyRQ9VtSHYBSDiSYa2i3Iv8Kg/RF0NjrNPF/kzBkWm1PCDqctbjPbuMOqWi
NgUNPfZNGZV9DKfZNXXISM3K5dzAQdL4FaGUl9NnMgT4PVzuR7h1VlEAG7DPD8bx
uRqLIj5E5rFRdqgMzvdxuB2Jn6nF/AeBkL5FL7BzSnn4UTsQnfB8hdZuvrHH0G3T
0Uyr7VSFmgul13hXryJlUeA966pvDkqll7dyjGi9RbtUd9ihZ/m03OVSPZwu7cc+
LJ+8mtd17L6r8ofz2Mv3BocHtqSBcoettj6Ud3YmLG7AEMonvLC9w4VCYWQZS6JR
DnV7S7i2azhbo/jUTzqhKbMTpZtXto37ebygGZL9APA8y6FqKpi790CgKJSsBSMS
Ib+U64gf55RdvF9ilQnJtcX3qnehVjDbwAYV6LoWFUBxKfl+YWshlY3fHtMdQXkn
xYzw+ErOXSEjwrYKcwHuDTAMGqNI1kywoF9p1vwe4l7Rvyz3fIN6QHmlc0nbJP0S
/+jxxsf6bNK06oBXkxQin5PtAeY6xndJRsCPufUbh5+CaiVrAjjESgP9HheuNtXj
MPHpw3QB7SS7YywoctjgUJnA2nUB/ny0vm04lw4iVBdOzAe5lTm1r0PDkgMXvEqR
bjaLNP/0TGUfqqDTdAtFKKQ1iesExkreAHXKdsw8iTCisWtCdVjI5Ezi9u2V9tAz
/awH8CuK7rEb1Y28rUquFMmMuzT3vcKep2ofC/C5SORHmpt9aIoYCZJVTuqWABiF
p2KIlwGVnDvi6WNIVPUlk+NCUf6iOMbhn7JhVH8/WeWz9EJvsWYhBOB0Doj23rMb
dJycG+tkCu5noI9bR8/eiisID65FTL5e3r1eEF/YtMtGrM6uQzsMgYgovOg10L3g
zosNCet5Vbo7UPFXxjT6AgN9LZDWheeyYSZMsMfpSU31tOoNzAakdBeqa8ya/Wrk
Ns9wFBOLvdBrjr92s+9io8raqUa7VoE4K4coyv2kgLQdIXDppde2OD/yqCnZKK0e
METXql75LZILOtDk0plePFgHUE0ifgpJThEBE02u37O1uZX9YgPwnwZ62r/R8akX
hHKoVtv8SfPMg/6tFUpi9jJ4LrC/WuQXFhzpDaCCcm58s1HiEr6IneVpRAiukH5l
W3wb5v2KuhwLO5VP5TcQXb/CSt/KWR9WpN0Khti1ABnBDnjxjvQIccMbIwwZOYnM
ME+bZnyRkqV1ATtaOfdufZ4m8dLtLrLp4OvlevKfY6rmtkUPTObl9IVGfhP6CYQP
tgBgl6iRlmoBJDNRzPFfHJhM4+LEqHI0fujZKiTnuiUcPEf5vlvtWDIZWEmv2qMm
2Z5GBigSoC1mabFLrNYsirNL497e52HzqvAkRy/ckrNXW9hQm6aX9sJ+in3HELvR
k+9EPwT1APUyyWhR6ktBtq/ROU/B4HDYQ+CEEucmVEJC1RZdC4FqEtRGOVb5onUH
19dquyF+JYUNwdXxi7SWSylNrsH+aYZJhruuIGjByyjxwkKFuwVnTpOqkksHDvm2
yyz80oQzO5rph46op8OgGegTrhBM3tU8/mR47bwXdteyZx5tQCB9Oxvvrq2fVo6U
UsEVAoNHJP+1+8X7l59gialcChgXM9/gLg1Bm/5/F7tF7vT024WHE4ojwKhcedYQ
c9qPYMaxDdO3BxcXE98q9dw/Chove+TE1sIUzIq37wGW7KTEp63BHl2/lGGLxIzJ
T3rmFCSqC6mqJXaSGHQdfNZXEXTdyZklpIpMazm3ucZ4aA1Btul5nCNui0LEnlgf
Egpp6f3bRqR4X/mbU+9FJmrbDsxjC2Zi1aJTsffmnYm/5aLSv9A7OHV/E2piEWSK
VIfQ525bGfQ9Ep25CR06fACuYZOO7ZGIlZBJwUNVQ+WpTQX4/JlaKk5CzzgJI5i9
vMIvLc0Z/1luWHz09frLkSzfjoVCWFAhESmssLVSw9LhciTPPRrwPeCPNTSVhz0h
ttHtUN1tsU1pkxjPCW1tBN6kXtWL1JgwLOtu7WeEpANQDGfRmotbJ+747KEC1J+n
ZsjOiLfXpejASDitcDEtwqcrl3Hmr5OJoQcE1biBIYr6Nq0JXSzK58MNNsxxyk4x
G0WkqIONTkoPrkT/uhzUZFn3QAZaN3Gl7nvxFVVcGIiiZkrS6Vkka93CIwUexa16
a+51EHu9tsAAN712HybPiekztChZuV+tHWvZ2AdCYXHv4IimAXY+XKkrZWDbBGe9
FMtSOu4J+8kEm7br/fr155popR2eMugJdX6LSku1utgWoYyxTyc40wjvbL+ZzbpS
oKwsWbVYsHIJa4AajZ2NShanRmyByKHT443DxucWMJH7jGAtzzEQBly8CxKIWMjR
vLiu0DmKr+ZFEdztjr+80HHtxaMfyc6rAyazU5THHbXl07R7A3RrKD+UHZaEXy4v
HK/Ebo2kLduOTLcAzx3smgaMlkWI/H0/SN0Qc1x1qD72QEmiNYRWmUKcf/nayRCG
FZsXycdqlEBiUNU+s0XvUrV7NmFKUWIa6JC2pYGK9FOXYggWFnuo2DQJ3mOxf8VZ
D3CmH2xN17QFL9vxGeFp+uLxSRgNlJa4f6kkSXBqR8Luuy0zf6edybCG+UEkr+FN
r3Z64JbsxRIy+PRO4Hy7am1teMVLye7ngn5u90gtlvG62Jpxz9n19vF98QRrfvjy
7k8B1BrwwgukRPIDJVZ+8WcERK6M9HfG+1YB6wE2koWiB3SQm0ADyKttidVyrCGv
zfmyICenn8n3HgWye0snxeR9TLk4DRY0OC0mgBNEAp3Ofnt6j9VnbUHosWjnzBrL
9qI/jzrQCw0PXEco3B2g+tYY+QCTfS8yVbaBPf7/Im12noA1hqRcrAIotDYapczQ
OFiO6inzOrXItA5jFq5Y2v3pMoI2qanzd3X/By3Ntad3X6oXe7iyjFI9/bjVvhg8
r1LcFyfgQgqmVvaBwBbukIPoITS5XCQzfMHtyutKB1fZM0cHt0ByrtBRqcR004h7
/N8yvH3Ta6Aie+411HNoCazafBJZdtxQ5nV4H89CV8KJABL2nv5btX58wCl2Ca0c
LaazY6gDwEprrw4S/YlqMCjXJOPMcLx7JT9Q1kHRbMu+D6W7yCXmpJqwhbtwXnrn
TsxcMxQwWQHXoT2E+d6k6PxbdS8Vs6QbrwxgMIFYASsnb7br2aLMY2VhSmUZOazN
Zt4ncpvVeWUl5z/AZodogpfFaooIQLbS0LUPrDTT0tqKHMJM38Pj3cGmMNLAMgCO
jgoGWHj3uhQH8AAo+ezsElZ25OFzCAqUzol0a89Yk9jn35EXp7ZxlCsAW7HhP9iR
1HoXgqDdZanZ3HmPthPdbPUxJh5W1GZzMavrBiWiS77DD1UDTg4olNLWTzqXBvnJ
PyOMosi6DOb6oVoU4buoT5mZ62/RkgpBUQVae2JoZKGIvAdN0mJTtQS2Irn/payY
fbL+Ot0qxyuPPwmGwFbETwnHS5jCOjDNrQpPwThm8GsWdbJagNHrjpRtkajqBqQ5
qiOS6sVhOsdAvD+oCNMFdwY2u2NY8o9q6g+69RDOitj1lN2xMxCBqHsuDE44Sgrp
lBoFBA24M8AlfRcbjfT4psPS61+V86X7cfxwqBhsXTDKPfF1k6V+9Q48WJMIMMgy
AhVgd9TiaJppZglpMwgCj9RULLc1oqj7GXQtgR130vSepTRQ+OnWVTvGRSI+96E/
RFARpdUnL1rQv3GGctaxxt2t4mL1PNJigq7XdoNj9/bM56i3ADxxtcGCXDuWCYWe
rQPm4fdlltfMaNF/8apaghET5no7gAfh0br8jEO/qjEbaTRFe/7Fu7H9In2bxoii
AloF+ncJmnxAId1kEPm7RfSCO8ZIjWkWvqv5H2jL4C+TzbHG+9iJYuEu1e0TnC3P
UMA7qe4S7YB4ldLgk9yePC8ZtrIChfx6kXzBUxluvNwtLPqGm6mQ9u3Bh8dw2Z/F
fd8ArCnr+iA+BCSEs8U48HpsTf+Y8FphLDs8E2YwMJUhjUWr2KZNx9ELSkeBBkFS
zks5G8jxOa24XbP0KV0hvroUTKHaWeshNiMilgfRCx7/JIK/zdOyzJXsvhndQ3L2
KX3km+bATy6bNRjhcnhlFdodo3FZ55AKXeOvQNx/uhYyBIxpUVwPxRzKVUENpK/D
8ColbXXsLY2JeBbAgF5W0CBsF1GK3wmVbgUSA7rTDav/Y1MliQBcKRrvK1ijZWiJ
RmX8OA1dmhya2Crb7SFXBP8JVhe1Ag6jfQtJLItjNavLbbjVVdzw+N3RPLyQdKZ3
jzHtSRLGXIUsGD8d7vWKY+ZPjMjNS51o+pwK+D7uuCIaQmJAjFLAh0xNNFCa2ie6
KeBwMckjWdAQwXhBJFtZke7GGfctIUZ690NAPbEqL8I/AeqgZxDf+woarxraCiJD
Sj9fVYYETL5kB2p9kSknWFsxmkZHsJ1VVok/7CvmvICx0NRnEgwA6P1mUuxCtW6h
X0nZpGHQnr4/kUhss6ic+yY08aOu0ee7b2OrHVPzIZVuWjtKOqJLRFmDbQDTTusA
uf9Sz+Xl3CDfU/orxmnJLwAnR/WcHwG9NNBMV3gNkVFqTEIZH9O7mBNJ4SXaGD/S
PdgduXFcqN79jqkM/WLOrKs6lKGRyIfZa/ns808PwRU+NsMZCm4SWuTmyi17Yx4I
AEISBq0D929Y1RW64wlM+l7vgrmS0kiQrCV5wIurou8kx567HI+Y9fkjdwmRK4ky
7JsndvUBxi6dG8U7c8wAwenkYHLbm79B3VDG2i7rPJHDQFJIuMfwuRvkJRQP9Fae
72hreBf/0eop/08Zj2DI0k1GOAH36eyseLeFrM9T5SvQpBjSvUpoArpfuuLQ4vS2
3t+95URG0VKrb9tCn+M2ETxVL00JYq6Ljybdq5sFwCliumGFPbSRpWWMBDCDsUTh
9uzbDvKw/etO7HZp296Ljxxjo2u9x8Z5I06v6KnDtO4G0a6r1SBlumPyVgKQMLoh
9ZkeMwWLI/gFbYYgp2zBFo+so2tog6bDHOrXVAH+oC8HuJnXvTpFZxdHbh5WCyQg
USmMGEAN9yFevIAnouiK5NyyjibhBZeXicglAY9kqtQP5bPtjZT9Bl77T7HEM4Ig
dIjqjCYW33Joi/nRj39vVwq9bu0S7ddueASvV9SLKXbKfa/lW9TyBbKvrYZRXSi1
vPxPS2ag4CaTwGwRSdE97oC5VrcvNyckHsMy3rYdRNzjJWxkdekht/ur3vXNyFYc
uDhkeCd3vx5fc/1wsUah/a1nWy6Bb2GCgKTWUO4qZOMzP5SLwQ19o9Ile0MqY/tL
KmYCDfoR2+ZPdWHngcWbWlYftdXWvoLxsPy5+pkjocqNH+rZ0oW1k11BHaRmJr97
iarslb+z1y8YHb6t/ZQcxdnJLO4X+A/HoJTLt/ADrro/D/P9LuftkobZ1s5kSZJt
C8NbQS+b9VE7kLGsjQ6Xhv3E0/rd5VGlmJuh/RDhWP7FcyZiAGhg/hv0K2ERS9CH
K8M6I6k5988eykUakbsDAF8OkXcLFrIivHlU9CbHlGFvQFtPcyH9LUkstuCybpP0
g4HJqlgSHWoidm2pocFgT3otEjcn44ZmrE/47Glb13pbp6TM8buaQAmJC+91YQYH
TZZDmfB2800hd3qNnBTmXHE4J2oJ6PqOojPdHOjL+lvEXvrWdU9Ev3iYqBdMZyne
8L2ouIi/MnOF8R286t5FiBV7/OAc+m0aW5HtTkyaHhcTmhJzUMA/1gYvHyZnJwwN
ANzTlLKAhc6OKaOR4GVp8rtos/F6ZslghhGR+2D8fztP4gRTodiyVf/QsVPB0k5o
hSAKlYRJBmC1tOcLoRMUMZv1EDoWr92nIGGQQGljTTx9TuL2zpkcLSkDA1HFWOOl
H/MXaE8CPsImXAPBehvnDpqJgZTWRgXj7jKBFqe37dpSoC3sm/etvw/AxEiw2nSx
gMB37AzJVfvNgm7QTWI7d/OH02MjVqO4ilKwWD4Ks9T0hPDB5VbsCms0cl5+GBo/
2K2kVIQoev0L5n+0Psw3cd6PIiczcv3g/Y4XPA74JiUidL8vHFSMwgBeQgxnYwQ8
KYfeY/RgyYxu92N2qMBfvwv2vLOEo/DE6vWQBBzKdAL60K/WR7QDNSioPFUaxHuC
+kY3LNL/kYg5Bo4OV+mKdUF/iHPRWgPdVKeZok9NdFwn1lINNOE/BmN4gysxGdcJ
wLsFdRtNgQDZgddiQfK7VN/tsYm4JlA7ZKjKeSPpM/gSwPmqlciX8Cb5YxqMtr3c
pM/anosHOLs49MBzoTPe44Et1w9McxbC95drOZUNHwiCEtmzzQBtIO9ZQWUm7zJW
+E7QSXPf0vgPKH1g2sZm31ZDBh3f8GbaYCXe4tqFfd7awwiobK3ia6ja1B+5qj8p
pW1JHusb/w+od9k4pq5Lc6NvcHc2rs/IOb+YFTZm0UN5OGDi/k4mMSUUl7Auo61t
tTAYV5NHvLshP3L8/48jmBOEnnuymwjL0JXs5krgmO4OgZ5b7Cef/tsrtWSvS3/u
H5tKjRvSHGDVM1Kw5Xpnix6BbRQIcHBwZ8i9FR0iB6Okc7uriJ7ZMZOE/Ie2UyGo
lyHYqJUEn5wmn9yuOTqpw+CBcBzuQxCHinN2LtaEx4NckZt4VGl7q5TiAjgytI9l
zwb/RmFI9gHAzA6+supMv+q1VswO8vwb9vAgsMzYTIXEl/P0XgvyFbTl3hgOT57H
7PRgo1tnG5dTKZ6XAEh/XwzIiso/dDRAufORpId/8kIaHa/ulhiNW2nlD5PrnIUO
2bkzwLdAf9V7JStynvd4j0QGACe0O5vx+giZRvc0ggzBnyf262YbKKbxXy8qJlwE
934MGC1np/3ST58i9rg2ob8Ul2ntpeHV7FXZ40nlIQwhQ1Mfgnu16I3LVJLq0f91
MleK+Y5XpVppfVxJSd6XhrgwufhEnDfSAuDIQ+PB3CJXUcKt3cZ/N2tUKfWHG4rP
aT4zw5zxIHTPBjbsNEq9NonPKX6Lal2lnLK+sv6gQbyxlVHdr6T9R66Rks6aVf+U
ZWzes7hc0o0w+4IbDvOe2oUOwvvvwmPGexcbxzvFPhh992gF83MtocdrlCYM4rEJ
kmmfxCWZGntSgRpKAKAhoEBowxg03nv8zfouImDWm6O2gNFrQKzbjRRQOmhZw1ko
ZUuoNjl/Dn3Erthg2gRievBlgJItkUyRGwG+IPASFDAbjW52em+Dn/s2fq3B+uSa
Ue1L7THOkoUyaxprHDHM074Oq/YUMMjSm0mgNsxz49hGa2woD8Bg7buCMZdX3iqo
o88GZK2z6dBuvwL82C9mZts6aa40G5higwXMjH4B807wkAzoKwbOMMf76frHQRSh
1GzviIPRDO9J0b7RRcu7mEo+ZxZF4xbK4a/Pa023SxGssaVAMVTLsYi4z0rwXYRp
TNn4M3uFeobhiKnPN0AF6fBQkurWn1+rF6d9v/QUzIXcIsQRK2ycBkatFoc6vKte
uejg/ONQrAEtaIuxJQ1LDGwoEB2W+nR0YIyrBzhAIMpf+Rw8i3WqHE2bLzIJXvbr
9+0hT0rAspDFfyXQHj2E6cvx8o/wEbVroDmejGjaF6kFWK0CcDZiBkmEGICj8+fz
StCn0GpU+5ifj8fE5RnWkm5J2wDNr63lnNsSERx5jF6uMGcNPGjqsS0n5XwFXP3S
6oqdrjWP0GNV4k2H0EfnBChhqjjSFZI+hDtNegEm77gMMROgRIRbFpM2oApOjC18
NCqo4wRD3BgNe5vg5LsSS33JXvc0r8hxvG3LjIp+610jY9UeGQ6GPiSmU8ZU8Mmt
3i46BbHFn0FybF3r4yMS7Qm/NWPN7ZEEjlQJlSdBVzngP59rwxG9o+ao0ST+mHbW
GaaAZKXWXdEMYP019b7bZANDfL+GlAUfWnk9HM0s9gYw3h9Yvl2yO2fULshl4wHf
9IdeWH1c7JzfJDVq+4L6bbHklvMwmObrb3Bs6rsffkhnecAmTurYZIu9TeU2Ezjk
kTD8nsfM68xopCqs2nnWCTE2dn+577feiPueq5bfze8D03nGqJ0WfTc3Wk3e0Nxw
EK4jnI8hKYmNM2ns1CLDxVIrn8cOHg9kWRS7otN9fj8scnml4vt4wbB5JjjWbnQD
SjXHl+yErbZHa3oqDzVHBi5TFVnPVZ9JA/RGtNYSJT4v48s0png834AZci25tGZb
sf0zNZWUWFvthR9PJIwqlTW4eCPdg/rtb54NcbIaca3Vae8yFgcFFBCiBu1v1UVr
ouqzS5S4c1SxFmy31cXAOu8eEps60b/Q5DYl6r2TBhh5yEdNJUyTesIQh4uc5Zig
mKzwM8znpmA6xf61P5rxuIqvHHPOXj9aSyPOwGSr/lnuTVyIiGjl5xyXskPzMHaa
ZIomQQcID9N16K8qKo9XovK/H1WfL94rWy3XCBPEZE/tvAEYEtRIvOMr4Fkou/LN
gKXfOQuyTfoiTfRskm5JVemfF7lknsQErWtVJ0X40aBCBt2iBxAxicmNAFNXOsus
VEbpuJky9LFIqEEC+f872M+07wrnVYlicYZ/Bsz0jLiUnzXZXte7KOBpClyACCQm
3hEWgYNSdO06deGKhGy2rJr18tBIjhMZZfKDa7xplrmyZYnaMoMrTXAaA9dvJ+Og
3xRhPSZBWlAK0QRkAOkALWUcoaFPGAMrwzN15HYHOlXIBp7aOPDEblSnE2aiw77e
+M01Ro9azmCTpQW7euNUy2W70EkRBGiHhW9ByXw2X25bJFmg6E3SYvFXmFS24qW4
O6ks6DnG/ga9ypQOt0j0LLQBr9t2+y5Vfl06N+8ZLipSycEDRnJL0QSWGDBqVAYs
2DawwSf0pkjFnEPDFOcfNR8G+OuJAYnkJGuDSlcJSuda1TjHhq7iEJNTajFhg885
qe7gfYJDVxcP0CeEvBp4F6e9Dtyl0uYQlno4NfvHEKyD1Iid+FDr2MSZuef0Nr13
FcyQ52yvG3cUfT7kksrc+jJ8QHGbRGXIEX66C3gPWa7yeWc4l7gk7ti5C5gWg/1V
Wy2f6vgLB+MTjgPY3HIkevmI7ukWoWkGh48MalWFZcGbO9KXhzzEHafEXlXABWsA
MZErtBtZemrhUJAV8wz3030FfWjxgK2ENlJlDmo8P49C+UaIMpAApZA8ZKuxmvOE
+jqRLuE/l3VupdPP8/wc5E9dVRe97hXT0nVFXHtptPWVvqq1X7txRh/yA4Rf571p
Xjf2jjPERfhtgUQlJW9m3o62ixTS1r4+uAb+S6sXp4/+DO/n6atF5eY+z6D7RobL
7VS18OD3y0JaUOXsBj+wQ2x1KmcDcR0e98RH6/zJUhPpF5i9fI7seZayVRT1M+qq
9a4M/blgz3DsR5eZDsFDA9ReGpfaepPSVg6C3wEhO9rXsTKkDNQ/wtOcQq8OBZ1l
assBkhKBMiLbrWhm2LX9WAnryUISYoZK8WF6WyC4M/vLuhAQGmmvc7rcL/vx8kuM
BztXUPIebvE1x03QeiBL8ME10ZhyxZZ5L94xP317/p73FEpSdUiidROqBzJN86z3
ACv6OJpYU9lfsK0Av2J59aQorJwgYEG3QkOa8gCkT16+nakw0MRagpn5U25PFFNg
26tZXmO7jOj56Ns/sT7rj6T4k7DnDnePzZM3XJR+g1kdnVGSst82Fc7g76p29Dju
piLqNShMyXbFdS/5q58OUN/DrbJTvOt6QhBfHt7ElxjEyr+VJibrkFe1RTjZopn9
N/tN52kARhZm3GdwakL0FM89erVt/ZWc2UUev4HhIaFBvrhvigP69vPBGxt9tcYK
yYkTE8pfP9MwCnq0Qi/kNXzhWPB4x+cqgdsIYl6YoE9nZyzkNkjzchrL3SPy/rFL
pd76EXf0VROxaPqXoM9ZFQbBp+6K5tXJjn5On1llbMAX2EUlaCEXV/9/Wv7HZq+n
AWF5s49H1lBstvSZBj8X9neYnatH4RJhNoa3TGDGciWAC5Rbrypn7PuzYHO9iq+H
dvicKVum2WlNElhYlmgpO9qeDd6jgFQvtG6cxRPpT1aYDCoK7rRckXuUNOy/eYql
57KhkY8Fp/YDEuTUcpuKG3d7MuAfFxzofvqTxTT1Hxu8OuI3c/hyxupAazlSzePH
ezNET9YlkgZqQ3/3QNxIEmlq+CpckVYSKi7eo90apACN9vDzQqttagGXBjNCfxVK
FQFBg/gVngfnQM+H7PY4FrGBchfHuLXDgfYjqyhSQqYZIlkMcaee37TG5YEactwM
9mD8aOKhY9tqT5huqjg5CzWTDnGEja0/tBsAtFUGrh41BCbVMDTUdNcDsp1swJIW
8DEj/+p5hObkDy8k/tietgP4+S8haukd3z8nKwbhwBeVWAwHdASQ3Fxiv5rjyUg2
U3t52oKXNCR77Lo0DvYFtr5zdIoeMvPCmDbuBXVjByG4meTHizArg1+Et2lsX6sz
sMOW98eEocnqlc2g6wDtYyVtDcYCFL1kxUqv2yJOw8GkyiTsqvLtePbhtNqHT7Sx
MrqyfxEVLQKAxi4/yCcssrO2cMHZ4SoTJUCoU8ovgGmMwgRsc9wb/x96jIfOZSPa
lRGLsKA2hjc7nyJeFHgxrAjxIR+vWN4131RMmRq15uQJjMUS9mK7jqVQt20VTPY4
j6Klqq28vWOF9h6rLR8+KT69FVeMYXP60JD26T03VQ0ELOEvaQRW8triIF2pXQFg
pR+Cz/TsW0zj3UJsvq13rykDSGHOj+XfM5JLD3MUqfopLQMYzHVg7rDOy7oKBeMg
R+5YPgeIzCWSnOXyOXGGthAbZop3DmkDNnQdx/QEH40y+PzrH/l88T2Fm9GTMaG3
JcrZE3fNycbdCw3AVgMjMs4s6fBltcemkgQHouN3m35RCwCpc3e7HSyJ9gJdAiIk
2CMTugX8mAH5ElMZ+tMaSXZ2Bx/rs0IEGKMePnZ+EaQod5NKkNXAtUfuQOjgD2So
SfJQZE9x5DSD/Hr/wQzyWRBNE64H1u8UK6JSN/3hiW2kMp5jDKgT5N3DNxqQR1VW
eEBYLBUcAZXYA5O2gy/LfIAYsinl13IQyjLQnB4vJfBrTiRXMqLm8U/jovNdlpM1
0TUVgQGYhSvnbUXL4ltXUfmYKhrHYiBrKkSOz7lqHCP+61+wLlq6c1BjYxCZgV9o
Rl9T8q3CaIMMTDTb7/1fBAmXEzQMiDpUCR1lSweE3OWg0JJk53N16yVub/uXY/Gb
H5IoN5lrdFKlkKOU9k2mr4ghUTRR2s4wnIXVSl3RGQxlQDepYuWP6eQckSAQo6tz
JA0rbwxBPlHobzVMlgp0u5Hpg5gJ/qX4zVEqPEbo7s6xY8b0CPkQm603eEl3wvwx
J8gZiMbdIdpVq2Ng2boX6HyIL3Na5Gre8z1eEb9zbKMbaPi/zDQa9Xrx7F92uefU
D83viggZiKrNz3EQo22GzplbOgCcAVRzxCxO3gLkMC9BVI8dALLJVrJLTiARqfJV
kvmod4vSlM66GQ3RrfrW03LSamfvmHfLTToK03azSXuBtdjCLa5/LB/TrVw5lJZk
PXfeNmDdvb2u4Gp5Ax0umk70sM5xHW1ntzeTps6OJctNUQ18UgSbcqbWpC7nX0Cp
hUq0PhN6znWEiDrNGgbKI51lpVltanc69kokeAl2nNmWUTj9rM8LRWd1Zyhb5W31
CpOn9EQE97Y9AuzHC1z7i7TE5OZVFDKkXSWoDbDJDWliKBjI3zK+eaN1ATwrZS+X
WSWyx2wxOkL7fpbtW6R4hSjudarzMKjV7AIe3FLndTb84zSU99eNLb/jQ1I6caFY
s/HCXSd4gcqU1NJ2A4oiU/LUVdYV2QAUAYYzrldedbh19Wh1MPvd0Yri2QZoT+jM
dyWu2EKsL99YTjYvpdGpcggwwymPjUONeAr7Oj2DuRgFCELsMUoJnr7k9SQCHMAM
qFB+pl47+PXxQPfdal8+C1AHCicc5aXjvkk7xbQMTwZLvC3wDk4P+7osV5KIJ8PG
dLQep4mAHtbFp6MoEocWI80jGKQu4gE1jdcifk5OV2eIJUkk2siUibeBglK0VaFl
ojRczhs4Cfm/P3CRLLbrgONDIaqpPKTHg7tSzhClKKkRUnLmkZIJaOFax+4OwiSh
f+qFm/iyVuAoarUCelxHNQWvyy0De1/1ZJH5sXen2b+0nXl1QPRoFBLkAljttIdE
WTt5QxG7N6hVsx8OCoSzmPxMFHM0LYcUJTUx6a9DU7yVtUInLn5q2XF5IMwITEfZ
FL4NWF01UO7ZSFCt/+x3NjIjaS5o4iAycY2PvWuc+etu6QYj7v71E1LVNlXZ69sZ
9JzmAaKcfZ7ppc9vACY3py/HUCNvzjLFbG7HYcniDTHlMUuk2nzqvLX5jtaywUEL
S4iLJtQiiE10LC1O23EzFyB9p4TkcADn60KqSjBzIs2wEMgI29p2OO+VX5VZ+oyN
uZx1c654hiwMS8Zlf384voawSymEORLFJDNAP5bNFstNFx6i6RHsSCycVe4Kf2Ka
zbbiwg+Kriru/uRwccLxWxqbs/9bZzLL+hNfl7FnKze1RkoLRFj/U22lir4UA/xs
Rr9JyjCsA1TE8OaNwpRJTnLPmTwRZhQcW7vc94V6mSpHGIAqXMdBH8LCHkrIw1+R
+KQ63kAa10ut9gHdIBRuLNLQ6p+6vO7QCP3+HHP0A0j64KOfi9/YChAQcQjd0IzZ
O3dW3drxEvMTXUCKhtBiBxzxBnU2QQSDqhLCoy3ZvPA58GG74hfPE0VcZFVxT6tf
B8ecjmW5h3O6pRxCmxQWTBy78MbT1Ibd4rW+ZTZKXbLQvA3KV/QEGTIEHv9kjXxX
/7LfZ12o4rq/PPXahOhFH41M83WNf5DPE4NrMe4Cfsg+rPkZzbEdyTZyubU7RuPc
AdD1BANqc5AUK7PuU8BWsRwG+NmMD9u6nXz5d9Vt9SJB7qH8dJODIK24vigwkvnz
I06jI00bk06GzGcsFIrtaTEVHUHE7rS1O3faNPs34/kDKZ6UVwqVN4uDZpLqvSvW
Og0Ao4OTo41DWYgXe5hOnJs8EJt/E/dcsNSY3iV+KrDNzbgKPYnsgrLbzwy9D9ma
XRJcvOa3Gd44iFdCV2oEk+n652S+r54FObpln+P3IeUtfDkg8b8tIbvFbWf5b9V+
08xLuDYHa1M/urpP3VcG7v6FbcDfVHb4bwLdPv/K3ru4MxN2BEBZxVphjM9iy53C
XE/GLp8NJy0Na8+b4b4duFiUBk0V8G4cCHYBsaGvg3vmh39fz82r80ldSU/OoiTW
nMNzA4+ASrHeOxxv+OEdSaUPMdhKOV4dG4Bnn9KQtTTmi3Hca/MvICdMQTvOhSaY
VU/DWT2DuYlv/LXFxjOmTl768XetZOGmrJ0co/eKWnKGNmpOnPs9KHsk9L0rbd5a
NKzo/7VdfxxY9Amw7mE04zWaiNJXkun47XgDwzgzGhAbTIXs5UGlJhA8QVe/LcGT
Td/y5EdYglJqM/NOj0o1v7/WTkEE+u1iYoKszJYWKNHiiJW0ZTOu1QiZygi99fOv
FULtpcRacuGJ9kZozuH4r5EHgibXjxdxqnZWdp2DpTBQJ/Mjfhf4WIg+oRAq1goJ
KIjtj3fEGBYAEJX8YFSU/Aw8/WFfKYoQ12gxZKYdtbFJoweuO4NAjQDBxJM3o2oJ
dCr+sNb57CYf25STdafa788S6K8mjDQf2ofj5d6/NjqLwdYhcFXBKymzBaKmj3jf
IJR87pCLyaTOD2kqgHdsd4ZHK/0q77fevVwRqFR1SAJMBWmENoDbOz1O5PcFuuCT
UTUVN8Tz1ABpt7wxhtyx4x1hsFCLR1T4SBGHigP3VJTHeYO1mjDquRg+AZ4HUEyr
y5N18j2NBVePg5cn1naC2ciVW5jw3HTbzBMFyvWfme1SXRQGdhawYf64Ex8TzrMM
TURaykHPcUdY6L9oBK0d7xgUeT4xTCeS/n8fD3/Aq/qr3JJ/xOMAV3cdum/0Hjfy
fqDHowsluy1kSEHuCP0QJ4693li5yMU9VyRD0yhMcEHqeOqdT1jsLggOnqv3hc3N
2hUnvyQ7r2wUIOl4pVjfW3TpqIhH1pUaiucEczqashR98ADvNbI1+ni1fUPpgoeU
/LanX2bS47d0kRB1+95WHclNIdh0RN7hqWjjIAuEvzwnFOgvIgHeX3hzTzLycVZr
Y4HSKd6VzPMhtdWY7He3WAehG9kV4aJOSYH8fj+VaDxpvpw1P/Np+6Q/UkmtR7t4
WZNCzbwbePxWo1sev5wljmFrnyrsfEB/Ozl9UWTKkAKCGKJwAp5FeNu3xK1sLexb
WMMGLWDAoiY3GSTsKidoKYzv3dVIMSUitglV6le1mTVEoPO7RZRehGkPagHnW4Uv
TJ9leJR6kJOG3rxoopcokLzR2LY8IFkePpx0+gXmk6JmHojyhn3EDMzzl5M2cNsP
eiZ9vQ5wms+tJezwC8WneAnUycBwL8TKX0SbXImcbqRD6s5bOsqJvn86uLcHwLGE
mSvhAIM8sUGo5OQJ5aUBvlHA4gvxC9Av5hrAtlAmfIMinzCoQPsU+vbLOvUpzeY9
ODZ1lgJf+g+8rsu3UW5FxNnHkquGaIKC79qQ5n/8xv5BOOgoPMJ3HH6VpigWMuS2
dvn37fmw7W5rpQ65ijNzfGjtgYBTVLC9G/nHVykZO9XNNmEz24K15F/YI6CwTz9A
JTNPA2xr23wwareyJh4JvyMtAOMWouUrVFoMDi2H7YW/leFjFLeDv0QdVQ0e2aP5
zFkoiJuuy/97/jFwskgZCSD/kdFQlDhYGyWZsPhneFfcO0h9JO8Ux6v5Dv7yBtEF
6TjRjFrDoRlsBBSf3yvx3aEdoyNHXpBjbsX4MIkBcRRsEIEWc7DNUuIxIaiiDprw
PG3ZMo4H61SBitfh7JaA2SZg4MYLnStI2kdnGbOBv6zfdUBwRXF/iXQHJBDJ99C0
aI5kn9aiLX31zQegJouseLVcYioP4ZrOEeu9zQ7qspieil0vApa+1bGtt3z+jT4N
WefU+SymylSmkR5E0mnH2QzoS14VnyeBdRsg4zOTheI+E9uy/fCnGId7niqUusy4
cOnr9QDTSkr0GBvRrrV53quMff0ZUGaBaHVUjsivYIUHV+JG+COPehqsS1LyyHUp
uiVleQpvvh+pRZKoSLw4esmJjTQK8nudWiFVRnfsb6Ta769H1V3aJIWvcjPGsjUI
mEqXJPAdoBnX4dInYIOtwCSfJ3yo39Yhosbz/gaXAJs18I+DyC3ttP5C0vYDkCoq
4Wl5ugI43t/2YOq8dmbFCL8Xz9iU1VSd4IY9WxfT1JMsQigPrbWTyeCS58jgkNv+
3iOXefyIjoDRlLP5tqV0TfFRGKpoxQKUlp/FEXp2nhu+NZXJ0La/RsIdlwBmsOtB
mHXPXgeHcHWP11sf89d1YIHa3EWPk1nOQc1kbjKezl6TpOyarCs04kFyFHfYiNyy
UNY4ocWzFe9T9ae+FOIvoMS5lsApj+mK2z80Sc/w+ZCcwtGyCvAMB0V0ckOVbutl
KK49SKVPUBeKRl+XZlmxe6Wo4zsR5bPFegL2RyRaASBODF2odiVjdCKF+2TDCiJF
2lQOlr4+ReppWbukN1INdeOAPjEwrRRYII2h1svjHz4wjkJC/F47Iayqxvya8pGQ
I1FXR/ZUlivDGurOx6jlcCX3vYuS4BNq9B8ko6G+MsXDqtTTfLyKubjuUKhNUtBd
Bjh8n4lcAD4cWk0gw2kGjWwhZB6MpFkTH9sQV1AZOBVLqOWLZfx/9Ix3L0Htvf0s
yr4lPD67CWyNyt5a3IAdHJLSpDk7UZZPiWJyZVFYdnIPonmdXRaAMfWGZQeT5jT/
j5+69N8o55ud3410qsyvHOdia/TraKcCbhb2sFeaqClrF+SqHV8Uk82NvQA/vGn+
AaLRBPSWFwUoBQJxNv238tQvv3ER3p6NGeZ9MKJdlEOCtTE5Pkzl/DnfB61HfOHy
/4XQv/EIoOn2MV5PuC2YVIS8YrZ8KhQH5dCwvPLd5cXqfSAfiz1gfCsBje+tZDrn
fJWUUy5Hk2FYkDiiLZq9Kf5/OtJAkrV3K0l9cIdSwqo26ArB6xp3xylT6Mr3d9XW
D2HGeZBYzyWvJ4FksYvij498Jw7mfxnpPNIoYa/WaTtQg7yKtOSd9GJX3i4vIP9c
RExGWkj2kjjdjj7lITvPxMtUDKHDglnzzdUI5BUaae1+gDrKDPpqOXjL4WkM3NIT
rzD86c4/3CozGZLUEYM7T/Dkn71fPaN2YXPGgSKhwd5IH/Y/L/ddHCMcWx1/Qc3F
GJB+1S9X/w2/bX5aif7RUcicWZ5fEP7UWVSvY9ktp8FvT5JTEOyJHznqVuaCQfWr
OKRZ8z1ZNNQPBaqav+uJcu/Ma9dWonCJ5ojyJRLajKRydD54Qq+JqhtCYY5ofaaW
ATnxLomEmB/jMM6nMvCpTZoFM3JgHOtg/XA13nnqPnx49Xy2hCAlKqP0wNHMISO1
/qGIejxov8M36byBTMpkPkahl6vTeV/AVvt3jI2HfwZJqB8wWnCe/8ef0Dn0LOLf
nfpKYTSlIIZzR4hyooC5pmTh8TiXo4O6aS2Yh1SSh5aLXArhjLWf1Ne6M5Qnyozh
w7hpQU9offKohdRSJJhRaYjCZHrIfsPDUlgHLpkrl9mGvH2t+YrCBTNK7aIz6ytj
RapD11cnB963q9FXImxPPOkKhgHiaU4gEV/Pnm+6Uk7qFRc4ep6U54fRRWuzXiyW
yXCYx+ZI4X4quy80W0CzggPKbzTJZu1kjYDKqI0Af65n1/9hMHnJ7uAIWohlug1c
whvJEqw/IR424m5VJbaK7qr4ZW/rKbPK5YQ3INrmy7m8T5IL0V72VxDQccnPxJdP
cTV/nGDdiZ3roG2E7IPqbwrq7kNRr1ByZML5RBpPE+6H1Y/bUhUO/XC+KrVglXBY
t0LTCphrTEjnO7S8hQkvaw9PxulUKnLDEiE0nk4LTXwxz1BL8HIaKzvnxejrMrOY
7zp/hKHH+Ksf4K8bGYM6hjMj4e+hrHkrXYNzuF8iRJ9bFlO3d8gAO1eOWN29uPLF
b0mQ2w4yTHEf4uHmRd0M8M8kG++yTiAdCsqw6CXb+BvudllujV+CpYqC1AeQOr+K
3i5JEb9UpQjnDgMLX6uCn4Ew9RgCxNadsVeFYxbAXihTs/wEMLbQWEr6G+eaD6gt
Q47+nshE2ufDJZYmme1/MmDGkCU9Vfh4BvWh6Pz3zAI/cPF9c8rC36fidiabLqyZ
+HlYA+ik2LVyVdDjzAWWkyZ1MGMrXnBTrmREY0due8JsAiQI6GhOQOi48p/fYrQ+
37sJFAnkZxbEUrc9omvL/vlxqetIwNOjOj4AclROZH49VhjG3jlDL3xnWGGvVaGq
VV3/u5T21F9KWlZQrt3gRVoBhZagllBHm0aicmHYwb1C/yAGcy8NoEhztfmg5mn0
5ozck25RjFVchgQIwMlYHHa256UUc9zUqrnpAZ/53NkgXHY/no55V9A6QtdHTVt7
L+3Vi9n7kguMc+WGxavyU9XCT/v1X1PrqxN/EBs/GX6UFsLxi9G9oIIzC9h5siMj
GOeLbZYlS939j69N11b01HfES1ELRtipkuE4ltLIq9haZnGQvBORPMpMhw5I1eoC
JPkk8/2n8MQjLhzXR1zMcyFRDGAqRWt3nLe/ALiU1P839VRsRO8Y+xMxE8YcDhLA
ioXBSwZNiwDpemg68XvLaXCFZRhQlaMfT5RvhSePHCf1c+P+uqaiAnC6me5i/L1w
xJeVu172McvA/AIqf+tf0uZsZ9JG4frx6f9SMt2VN66NWLJDxfZkDKnVGGe2zI2H
BiFK+BJBGYrsJ6QtNzSjvHQ+VZjUE/B8HlMvInaMKVgrbgCoTo6PkNXOikwR8tVe
XBexc1xYc9bUCpdUpiTnvsaz/RgwKi6cF26pDeBMdpnpXw188dm2k9HHIy0fjVUh
mR40bSO2/Lnwbge1SKIc4oI5XASYkFlP/0YW49yom20U499P4nMNcIGioZlm/LRx
gLbbm4RlRvEvGl3ymu44wnScrdFL0oD4PSn7mIv06AvDRpn/FfER3SaftjuHzK4S
mNlc2LOX6H9AUBr+APARy3upcmPqYY3wFjXR8lNsbP7/mprpYu8I1NOexdbZtVCe
k1DyPCIYaWR/AYbLSIgXb2z7tceXSwJj4RRylT8wB7uiEHLYgCqpZHsvb+YwDGPf
YRkMcbcsl3GVPKHqPv/RaNFoAKLZC4C0P4gj4GTWlS3ZsUQsarIWjwVZmiwXDwtD
tJxz4s5UNnGTc7Xpb2jFYuNdGZOGkzDCJb9imRP7eM9/9LPLaeZVbYrmBf3X5L1N
7suUcYJ3AgcbUeV3yYNsvRqTiFb9Lr600jfiA3zPKnRmtRN6F2947KGH0LKTWoaF
uJNujfmhRJxiO5T4VNY9T2AEHrCqCvvRxV0DVWkOdsWX0wJwELJNsqRziop80pDc
+u9sOpeQj2+i2t8yzb1PX03rj69wNpOVKqRf6QFXzY3JgyNAiRq4y6PBVn0yFN7q
/xbYU4V4J9pR6p9xESHP9CK+UA2GQpjsOv/uNejWgUFiMFuhf3oKVTl71atFWvqM
AQG60RKR0pen9CZZ9hjxcemKBAWvj1TfBpZ4LTnslWSkLou7jBaUKao4aLiBsw+E
3A70Nnj2yBEaZytFaJTutXtefrM5MTg5HOfYBq1Be8CCnJcfUYcBR1L8RE3kL4WI
9JzMJ+wEvhxyed7iipzY7uki+tjKQl6HzyupYop9h75aN+Fc15H+KhglXloL5BGc
WmH1O/p7uiz//pr/BvP14j1A6UYLR30xHiStPhvQT/0nlWZW7dHc73t9I9qw58CG
hjbEn2183FGy2sVESlUQKHnC3KHY0NHoYD+GSRCODlF/gg7zGkNRSZ041aRri4Vn
E+aKHBRufcyxIowdIaMgxU256GeS4nG8SRXEyXx2OVKFI2vd8i5y7ek4YEx3d7q7
1gwWyjYGmWu77sMi4hF6nkxEDnd1Ms0YKBq9sOpNBtX0Dbpv7JNIu2OIuKF4Q0eY
BkVn2+71h3IAcAF4eYPNajNnLkyqZrH/e6+0JSEkOUlLFDGRaA8iokw8u7rkHPmY
IT/wovp/Pl61AJgub+i+qOLHwWBZyrpDjHzvHLyv1rIGLoZwV5GR2cI1IVwGN+S1
L7R61kxoNp/5o38CLWXajmJH85NaDU22hgiy1VncFiGYuUFRL4UMEnR8OpU2X465
XjQdjUgxJOvQkcanrOmEW33r3iFT9VBy9oNwBk5jcX5dMa0mfEI+10Y3tLF8UE7s
zbRipDYdGrTEx2anVt1nDIl8ao0buXXJimmNzAQaUX/XltScN31mD5mI/9bWuuLG
ZWFyF28XkG0yZZEjg0RiReg3mbBONDOaJsmnBxLhGYGF3q6ShTuev4OYRTGSed90
WGXyDvSJbs1axwxB1vH8Jfi2HOKpaKVbxIbXGR8DfMVI/qanGLzOw2X+6SgMFl59
rWNWvt2MBQOQbhau1ipmxUzZ9xrbuuEViBIamJD95h2lUHDTZLkObKGyM7nxXlfB
3H6pddWF/LP1jzJ4Ya+jwouoxsAs72x/2OXN/Ial7lUaAbTWXAmMEg1UtUtrFBIG
wGxeQp183zSVdnt4uWAWv/94GSLeSoeAkAgGzgwHDQo/teCjEWX+KuFOtPElffFP
vHd0WaLmzoIPmRhjTE+lf/pY4irwsccp+iLceOFuJc2B9RiHBAPf2eznKMXEJNg+
R83GBG5QPA6Gy+HqnVfH6F/EMyJxGEyLaX4cA9Lyx77gRpm1WsZk/VdE0JlpsXhb
Sb49rIIz/PCp0Y9wHrFQq/nzp0wH5Jj2wSW2sytj7buqflgAtjIpFfc71LP6eidL
RBJZSJhqUmqCD0+VfhHz80tNTiS3g/FZCJVIYMunKFFyfLmX853HKkI+5ABlVPRz
z2Zh/M5blVEnksDMSfh2yIE/Q6eV9L+Tz2Nyg7m88r+QHke5kUTvw4fflTLWy3cD
WQqQKhj84LQXCw/R6gIGUONsBynqLXlK5WE8dazXlEbmYzG0xnUYvdUGSQfzQm94
tzZWZICdp0ZQmYcl2LfbfNOopnDI6rDVvPD5fz+2P0QZK3axBIabwNUbpXy4yZ3t
06s4z5tNNXoRJz8oYxXCxRiHbUzmxpjGRmGfO8TqBKUm4MdDn+Vu8RUg6s7rQLNa
H7Nji4i1BhQTa5PqzlTfvfhrWU9TKWeAmQ2xAn0sGWyDBhRfMauwtiJDSh5bJF1p
jJkRHS2xDsbxKXjFNqFuFb7E/pAAHAJXc6vPA5jXJZrbHoaAfON0AAUohl0RnzqJ
vhaDMzFjVQmDr50aW9wR/UAr32wdemYT380UGVC7u05hnsv+nslzuDv3ZW0yJSsZ
X7gcJ+O4Lackqx8/wAcm0ea0w+G48WFZjcHYB0dUsvpHye5oXTj8U5henkKO7nfo
ZrzHUeDd1b6cKfE19oW/9iSH4bUP9v0Mh7dLgzqU1qcF9KXOBnGhVdm3qNEAg7NY
Gy5sYuCQybHQhMcV1WLDGSjNOFWGfUF7UStiIm+sQfnV8zFaxUEWR4kYjIWZMMaH
/NAwusSyQNDuCWzS/p/k3xtIld9aBwxScmFejRPueUBBUeGFqkLdTUjkPeYVwpLG
TND9KlL+GtaVOiMSce9QZ/1vUkyNtXsl2DRBZ2AllNSrEwE0BnOSjOHyZSLN17W3
iCkve2vDVYmttI9+HHj5WJkw603C6xv7r8pXQ2vsopZ/9gKgF8G6RiroUwmQqdwk
qxFIG9u1vKMEJrFqJ/YYeN973ZaXN4vp2Ax+8kSApROZCRIXMvsNFOE7q+rtEZZo
/j5PR6OXqcVnOYItoTew5flKeoEGV48dCFVWzCjiVTnYCp1zi3etrS8U9VYi61U6
76YM188lc7flQIpAKnPXutFvXf0p3juy6A0tLRvHwehTG+ACQaZCfqV1njHOId73
fQqvuCRolvlCYDx4KUQtfbFem5CbXWKsNBzzCGVy1PspAA40ED0H5lJtBkk9nFNO
x9TJ8ZnD+Ro8dYv90uCX1+AIjw7yfe7Bzj0ViXdydHRTJHs/D2YttWt6Bf1L5Rfz
oVfam4aZgSc4SHNHih8tg1NYVkxf2xSmp0Jx034IgqoA0bKvjFR3ioQpaCwcEVo6
KEtXVD+IQGiuRRAhw7JSxHlZKZMrT+CnXPobMfWBipDkDpTtiASalmBPVGTJDLYu
ehSUSFKQJgaq+IWDyqgIAK7LXJO+JbO5RW78UW293gW/+o3SX0cVGiNoZlQmBbev
Quumwu5JP9IuIRPYKLu4AMvCrD/URYIXdIWFZEIvjFdi33cT7/PdBS0/sr5q9NF4
GMUjSZW8LVtP/QIdjyF+7OR43T2RXT1D6gkhncUYansOIONyoZL57IPRlPvKFHPQ
Z/Tj3XEuPzOee4xIV1T8g1gBTMTuhwZ0mDJglQncasb+VPMJdIzOH46j2cQHq2xn
bfyw5Ismeei5goGgvMLHtVOrYstOCzKPTLpb4Qfv4iVpO76cKMrkc9UKXBTkUDJ8
vtoqgeArAuHSdm0vd8bR7noeDa+7v+3r+eiehPVhUVf7kjiJ/QkQkS5FQmHD0kH/
425cWPB36B2WPutwwNfNwXkYNS4qmYSKRxpb1a1jAd/2WcYA4Id/XVJjJXt3etUJ
1zRr5UuV5BaKdRAn09T+CKRXd5JlB6g3eysZWXVnjAGJnMLAhKMZtv8sxRiG2poE
3cj0O2B8uzpUrSD4iitJDgeZi7SJwrlmbJv1Z96SjL/T/biWe0Ju0MVwCLeYQbOz
KRBJo+AVaPL3GiIHD593LGJvff5XvTno/m4kaV5XGgglbmX5NqVGBxHTeITuq/s/
+a/lRvbtSlauNLqcrTxbAiGkgAoQpFAMJezcWLC7EgVM0W1dMQLVn1snqRC3+Lbt
aEmzkc19XkMNEsSjWXMtnPLhFODl0NST9gDOaDZE25wIB5Lt3Hpts3WsPJslrsmd
oxvSVHfz9AeEYLUhDFYIiS76VyQcw2lwQx1S275Z2UtlRZg/G57O3I8iFapqfxA3
LFCQAKpeeQjfSy/RvHthkBR1o4aVoXIOiLghotPKmk3obfiGK3fKWSdTlMVsledT
+FdV9B/m0iooTSPv/RtZheMIu7NXmJSxDtHlAx8HHEEpjKyM/O3huYFC9A35Wucr
sUuHVq2I2pXjAMwI3ac20AJgZ+p4tBbGTZUKeu5rCT2e1kFLY8xDvvT6XPTFvDOz
f6rIc3FTAkaN6JYLZzLbBJKrCaR2Nm+Ml8qxH6Qnl4g0YfKriqSrMpMLGA/BdqPr
sS1XVq0V3iHfMiCb2AVRUO6BMhAV0eGymCeRt59ao5kylxs+Tr3oonXm3khVsxh4
z51GPAxQNDvpuOQH8YZX2jUyDpOWaoKkpcRHZjuBaaW6idPEIhWn5ay416ks8D/p
CfNsLKbmCDcZ+ECs+SI8Xo8kLeGqKJjRYmSYarB9Szcy7Brjdvfv8Gxfu7lopPxS
rE2UHDcqrchvnLLoevG/ek40ggfQaIWfUGR5nic/McZ6sTw7lu9Ro+8rC/dHssWL
8Tz5l1KRpq+bE+YMuoIJEa1RU0KvE3u5+QddrUW/jVMNIoeUPuHRCm+6Ynxz4I6v
ZZFHM4760l78AmfsMcaPZkz/hDmOPgs7tamA0dAlcRTVUM41HirBHppGWa/DFe7n
ElrIYjxF1U4wPVzFAlOPvL5k6hv8akw3H/J5Ua1i5Rpc0WxZTRPUKqfORMXSsqap
mPiNgkViI3njtY/QbbxxKqIDk0cR0BFkIo6Oos+AG2PZoSu1R2ixuyjGF602LITt
wQNG5C7gqIzb9tZIFBQWXywOhggq+oeDWCzv7and+HMy/bTFKTdUb5L+S8GAFRO1
Kdc5s9euPiWXA1tOawUCqrU9aKuyIqFJtv15fZJFKY7AczOMeog//7c1bytiCytP
dPLG8Kj6JALlWwI1gmb/K0qSe6JcMPWRGSLr8Xn4vGieobgIItTdBHi4EHQI4LbK
+B03thFBBnIDPgweQba6v5IE5wRl79s9Gyu+QXoUJQkKZOIAdj+dvLH7PsIkuQhC
PosMB/gYrhFKi0nkiBfUltmMqDf12fPNkmh1QaL8grU3PkLqmNe003mNX6SsxC5U
5wsBTGaaRy9iK62S+oRV+rPQXpAnzRZLY60gn7R406vKY2cDlzHZgpSxvIUgH1ry
era/Ft24oXrd+bDvHel7rIsaDO1R9b9sX4WRf69mNy3Tpnm0PvCkAOZNYUz9fy4t
5Fvr2UU/FKOsDCNu6xwYWRGBzFN7u3fDmCQMJ7ViauDpqTb/1qcZkHvjwynt8I5+
G1FqrEeZXyQv3OiqUfMjASDjlxqSmYcOuN4QTizc1i8juFl5OEXKsWjzO6SgbJsR
KrA6gSCOE+tmgf1tST6spS6XKIFmqqmrEZ2T9ZOilVEkwyuTue8IIqvpB3P409jb
bPXeat5OQxsqFKVm0X2auHQy1Z9rUF0UOvt7ovMIrn2z9v8hHHcywJY8uUux3Y4M
L8GJOZqe/qBvGFJ2tcPUac04l8QELldDkB56ukeo2wtTc/bIfJIemkvm53wWqS9h
CvZaDH/wzMsZH8JNTc3ENjCvWKFWhmqJ+iHosAUc/NfTl1noaqf8Cp6ii64ai8h4
mWsBZUGJPOI6hZFY/NV82wPpHlA3fmfypbEhc2fO2bfIZZG6t5g1XjtBeCuWsdH5
akZP2+afhOS4LAhTgrtZD0SaIXeKJ6G2QPnhRg8+3aR/Sy20v3mfN+v+FLWdMzDJ
gYJ98FveKd7w/ly/Ku8nGF+vIa4ieqFxF130ztTMC/47gO3JfeqxF6XIg84gI6//
IGUp9oiVHubA80HBMq09/qMlDMrok2ebObI8d1kAsTAux54Jpq84SRP7kZWBgQ+U
yAxYp0GczCw8f/PiNfJtgeRIEp/b7QHklZ7n2CVDw34aj3VkPRJD7yqAR83u6/yq
LM4Sm5AcmTFjoZK/tCA0altRKj1OkcUzlgOGdAF6ePANmorS0k1lK587Usep4Y8e
SifTuEJiZJrcuaKdYm/i8Psf9i7wxqDjOJmZcHMLRHgdlJ4C5WiYAXdtECZxqqKa
lxD9EO8xiO5JwHlj7WFlTUN+LLU9ahVhsLoeZ3FBBGdJPYy32xFnoGFnsLMSKzR9
AmqlPUXps7Cwi3Lkcl8rW5uQp7UaqiX1FnEcTt2cgUri2XkXS/kMe/bobmNs0job
NkbzOPazf0l3WAiV5qDJxzIsZNDRAYYHQIVFMcyC2r29HTtp3LC149k61oxi/3vC
PK2tRq83UNfUZ1zCDAuHzjtzdkRnGb/kbZP9G4MDUi47c4EO5lkgIWop5E2Od3LZ
/EYjcQibTTsdgOcQNeJqwTJAKNpH+hn2R8yNbsx25P15wLq8We1Nqnl7AhqSFtQL
TFQ9uXem3Vjge1pLZrnW+KBroJmn2lpU6rBKv6UhT6gVDBJgI1QJuOIAvHRcJNHX
JGmD21d4JkGafAE/ob1qvStA/+z/vS/iplcoUzU7f4LgyKKsH2HVc2POI4m3ep4j
WbfhbanAluQvY7j58Aa52/HvnoMStjfV/SZYaKL66cqrXcbV/2JYAZVd7075FqUE
KScZa2hChHrdUUZTT7EpSPlRYLOJ5d/Cs/LV+T5lYC2lJFvke+0ZL1qK5FgqJYqK
qxyIwLHf0Er5rUlzVECYZG9IYFPfxl3iB2+hst5GQVFt2JdSzyHQLOyUFT9K3m6t
8HKh8oc9VnrWE6DWhRE7yVBtDQFGZHbFJdTh2cJ7Cnoa0lN7m24UDdKfjPF3vU0H
h0YNKJL1nlVsWaCalEght10oQNVEddmeu+rmzHjIDpPLu8SIJmzkS6ldBAmdZWfy
0+DREfNimxOV9zt/qZuYnZef6GtZiQunoIu2dLzT+2A6Yrvny4Lj2Wev8+dl/Kp+
4EDxfOQb8Bsr06DDqVXzQiLf6bx1hYBe70gmxxdonXHDsZK0pAL5YURUY11ASbQq
70zo37mDXxKQFXSaURJ7hOx/zMTO/e82dAGus9+qT574EbCJ/hSkq9feEIf9o2tk
5FF8T3jm3fFSqlmK5PK4AexUy5CAulqBgSIUTGKDoj37zIhKTQOxbOC+ZrrxWlKM
JB6TeNOY+HeIz+mNknkqMxa8bR0hQwGJMvb2cX1DlNTuFB7mrAlw7vuMbFKM3lgY
kwUSVWjVOZ10eqPKUdz5hhBWzSqYpkmkHlorHRkqr+sF0SjZEh3sk9KaJt0PrUXA
hIylodHOMuP+Ins+ePjc/11ZzlaME5H1wQQU5KtcMKhCDm2gJ5M4/6rnEW/XD9JE
bre+U7K9EQCgIi2L94ZQHjaaJmIpPMFvzC4mDoPxT1LHUy8+zEjKhBJ0MVK4C7o1
bam25behXnH4KAi9MeRjO2QBJbPTWeu0Zgg8lozplKJX9QPAzPbcXfZO50kkSkRV
gXDDg45PfCXd8e/imwGyjMOMsOny47zg789kuHadh+6+eQQZeaIPp3QyhvMJmTJF
Xq0An49+P5dcyZZskpkAPLv4m8MBKiCKOpm4hLUDnm3UR44Z8+JDxCoOPQT8ZF6y
5jtBbg3iSqw2sfJHFPWgY7STY0ij3iTPw6A2DOK7K9gpDeCRp9/KQKGHq24kCon5
bHnQ3H7bu8xVzHgzSrk9eTpmhcsp8thFMvxM8ebA1gnu2QpLIUfM8a0WvDks8gYG
uE/JbihhVVLRzFjR3NTLcAyEMqN7fQsSv9URetHT03CNkRn+CmHt9VeAcYK8xZit
vdVWhnScipVafRFyDBGMqYmBldq760hTWyAO2lOxCePXzSpJEnQPHmedNtUoTbkq
ezbp9S2//9hjHVneavBva8w0buzInZFzJk+gX/CYgoMx7lAaA4pwqL9x3OHQg44l
bTsr6eU2S9IlmDQ6KRAUFnkuwBXoYEX1ADYD+9NS0p0Q7ztuUbxSPk4co8s6Rlyj
Wq7AxotLxFgkuys6lMIvKeOa+RMaYppYtqDNHBmV1HcXAzlap0c2GKJM1vCgywiw
3aHGhW0R/R6aKDPlz431JhY8aPYFaA5bjeZ+0zE8uotTG5ycl/Od1nJ56FgYille
pZPvIk1VL1nj6kTPTiKg5xDpS6YT08vpnYHw5EDHj1sbePXIITO1PC1YLwr9+tg4
nXWlLTLpZ/jdM4XVU5UaelNYVBWW66BuOxnsLkFKKhYIfE8gyyyleO/s5oEjCGGQ
yGx2X282YoAuQTHY+7RRieKiHIeFA+Zu5wCnBtITXqry+WPq123r2lqTUDP5SRrk
i2FpJ1hvszhBlD4vQ1ua+fWHMzJAWbLPUj0d1ibCkRc4YrksXyv8dcWiq6KT+wxI
MZdOSYoG+rG+6JcaH0FC0ZHhlFUECBO1bDFKEnSHW90Y7b2tRvxReeYRwpVe42m0
wWnJpnNgzKcXGP89YBXPIa59z0b1JoBVfzSyRl0cc2lFgRv9kKfhlmqlFzbOb1ZU
m+l/RMmH9DM/XHMa/OOvp4gY+lZ2EEdyC7rTW6DUuqoD6vErvX7RoJAlvOvKrul0
tJ9hycrCOKR2ZA9NpO+h2K0RXPcDmd/lqJAWNrBKN0/TWI1Yr1vYqpvsOwKuRs/V
Qs4Y5pC8/TLMIW4slwF/E+op+ctpbPtlBrWpLPuKwGhlVKLrRzxoR7usCiABArRS
b5PUYBdSjXKo4VApuNWLh1bDkUTWSivIHNXJeocvzG9YMmqtNKWb6njE2nV5UCk6
+QroB2dMphoBqC9Kr38f43rNsriKyONt/bSSZi0GzIx2GUDz8/2B2SEUcLDCvx4/
bqxZLvCaXGXtsOE1Be8PEMhbx+Z4JFRgLSe1gvi5j4nvSFGiPJB08NUVVCSKvQk2
ltBPW7mcHBtoccIx72MB4YJgpgEhod3SaTOIxW0pUVnkJjoVpFCAaImATbdOr3Qy
R1klo1fOCQqOKq98v/uAqf01yE4k2aXkgPodaKJJ9FywNoQkCnDS6z3Z8SQzRE94
s9n6GeR61FoD8WueMspMgUl96GI0T/bAJNmn34fKVHmpOOLOL2w/JJb4tnRy7+fW
9Zwwb6HLCvqp+f6X63/JGnuJzReH78TEJdmnMc2v6CTFhyNXpNlv8LA9HROOUjQ2
579DTDKOQXl7wdzd2DNin2LQDymqXdkr+03ETKxGTYpS3jCbYgtC/pSbyaUkakPw
movk2kS/ZGwZBaMDwS1+XZw00TeJoI6MrDJNQb9aoI+14GvL2IakgAgPV95nMHiy
OztbA3Oz+HFOravXIEj9HlyO6TxH0LLG83L2sEkwwDQJMeOKyRUiXTU0h13gD5Uf
C1d+qPAylp0EgAdK5Nb9sLd/ALwL6iDN0fYZ2lliosJWesSvwndLH8paON796f3n
skWWqi/C1NKuMsJ+AsjJ9bWz/mbhlVlV36S5tYTIp1iyC92iBl27MSUx+d2ox41b
7o3E5Hk8T+kP92H4GHG4ywgNQnXhj1+bpuqHo1BuAYBXGyqOER2lKyi3bydiMMsM
Nq6HdVvAIu37zULQHm2NgeqqzeshWwmAYQrxXGfnYV/DCNj4vy9FniM3tOjENhqh
rnq1ckTO4qaxwwib8UGn8vEUH4dzbt6Xc9d7JKyEWgcBWZJIV7C73bMFviGpfCxm
ipRqCLful8IonPtdT5ejK8AY4SzZvQAr4wTDT52gooeaefNxao/an0M8Izo6sRcB
CBpk741n5WAbkXSpnxmQz/LWEyUCfOdKb8zmraGNXZUm/TbMjlZnUWz7dSltJPCe
mi5D+f/RVQFKCbN1cfMrU4iUKsLvSTlpgRN4Nw2/D5it8XsV5meRtd+MggQUUy58
L0eF7OhGg7pXbd+uVYKQM93HCj/FRnUP2pevMhP0HdVW70XJBdymnwbepIMAftHm
crO1F/elnfjG6W8oYgCeBGy/LEh9E0AbgVI2hm3GXUiB6z55TJqZLb8a1FsQaCbw
LC7LdGGHYTZTyqJXNSBx+6nUnjUOgHFrvVBjiAjPHq57kilA/EBo+uTnHfjzU4x+
teEjof6/oxfFAU2jBOBHOTk2pbX/Z6IkO/6Cwe3Nn/7wbegFAI8g8uWMGy47F40k
UtDvbE40UClosHjSz9YP12Rhvtrun5psnCzKFatG8saeNc7VJ7nJ1SyvRMGt4diw
Bm2NcTWZ6QTFp4rePPLcdPDBgH5ebXs1HQfp2uVhL66ctc4uF6O72pcBCTrcbsOO
0uv9m5YCwl/fEHTDWxMu7G/3XFWSNDWV6LP6qG+grPY7fA9p7VUF4mr8TdI0YkV2
41ksZXvOT0GX/SEKQODCSuShWraReqbFjWUPhrd2Ic2MOImU0ml460BzLbDnuuIK
Clsewp3U2KPmkrDSWeh0MQl1swxFnJ1OSi4R5O6VvcMtKSa76vvkGiH54bJ6+qcT
v2xhn5aLOsx11/BMstvQootjOgmI6DIZWZKtcGUJkLQvJbvJVNo/gZrWX1VzJVRs
CXXEOteuwfo9hB6joZKmcmCBcuuWO6tJSpiLeaQeTKFpa5nH9DB03kASjQcxNso2
TbBC3/6V6RVJZd5h6PZIMuHRPKRLYm2X10EtUpPyJs1z7cS6CY2nd5YITSEPLAor
R1lYOjnSucX3BWAYQ2YMFmX6Cjcuba6n1d9sfLSvdIka8+WElWhVUHZNzoPw9zbH
89zL1PQ4mbrt2gkbkredk429/8tvxlsIXWCF2QoAwu8bWSV4yxRf5jnBljWh7hFY
Z+xYRjPA1APEFB7hsDH4hZlCd8iSioy0o8pxeWDiaXDEoT/HeJh4Wg/TeiAShFXN
j1jT8Euqp2gCHFRNsZYhzybtAy4QwuKfQFqNV0M+6mC2MB3ssRdtyCdB/RYltaNY
0kP1SI1s9WUgMgCqoRfkyGcSd6PRQXWmNEGKXYXgW8G3XpQIKg6tejfrSMWaM0BQ
N6vkkuHzqSIdOBpjkQe8bEkT0fRXET+MZL5656LCsKBz6VW7S8BZ75M6yWw+VPSB
VUx+o7JAXFWAqhKTFlvfiueieTfuMXiks2bDCNd2aNT//sBLVtv8k9oXKkwMafM2
yRP5+zoPxroNHJGPj5Xyf9ejMH7RFp59KXMOwx4CynruS/dEy0xwJzRMxUPmTaUN
IKCT8pv4T/vdidgmHSpG7YiGxc+0ysGgrgg21uzK/hRwZgaYpm04TNp9NPI/rU8r
/XBieG1u4vIelb9HtTYnAiIFV4wLgR2YkilfOHbbtYu37tE/6fxrkfKilc9t8QvS
xrYlXU/lbaBazaaYpneS48zQJySrZYxrkb3MNGDdvhstv1Ixd1TKmc3YZCKZj51B
7LmR3MxNTHYOuFjEOHACJ6q5if1zvaD21bX9LYlO4SpPzYvrqWDacUHOe0n1bMir
rqk/XDKIrDirB/NiVi/dOEHbUN53QOxnKHaIbdT9L2wFsd52crtC5phSns5ZPsrv
njfY5AE1YaMLU9T6eMIRD+tkmOTM+WFkM5PiAepOeRbT0R6gqoBJjrqkIXWr5+Sv
F9CSbSKomaLD//bapkxusW2olFTdBeR3ak8NRGoMjm3hNDue1rB3C95hUzSFvfYz
3Ip9MPA7tbTwlW4xfi+7psFYcfpMbbvTLKr/5XMOw4tCbFaKDRJHARsnW3nj0DxK
mW+XgmZQHPRbeQvfFydrbwD3lj3GBzsYJHNcqIFCVeCH2e7d5u5YXiIJmox+PaHh
jKHsNOZhAjyvt03kTe1LDiCu4k+WnCyAyEHBkZz5r+0E04z8hee7Ui1hmHeZWm1j
9/NsIwqYOwRvQ/NbAsEPbOVPypny5a+y/ee7H4yongeqaSfKnyBd0qZTcMnDtP9W
pwBoYpWdpzb+xdTHiWo5xdJ2zTSJfGUBvjX1NlCDIcReCpgW47Ss1031QZl32I6/
QbtCW0ugAxnSC+z0E+GIbM9GccRctYjHob5+eCUJ+gm9y6JhjLsxMmDP2Ri0/n80
qFfpeUVCPT8BCIKWE5+8EAZ+cAE5SoxD5vzmalyzThNWL6mSqJ2anTbIf7P+nF3p
BxBJ8d/YqLeRLowlxROEvetVIGfgFvDfY5aMdrzFjzgygzC1dF1LmOGv+UTgNawY
rmcbmnsGcYcXRimjzmPm7buMiFpfcBXVp2PlSNlrZTL8F90lxoyE1/CL/S+K+GOx
0udXjcrxYtv6Xd2mCxc1yryM9ejr9Tim5PTcuzvotaVhD4+VslJ17d8OXkME4vlD
5H2dsKnoV7a2mv8Hq3DBNFdbP/XhxtHPfD1JHsk/J1UoS8WjSAy6+4jjPePvBNGv
U3qN11GkFMvX31rRxoM+LPeYG6p4HYQYSPceVMaQut4X5df6IttPRKogof0TZxcf
b/F3/O/VEaKKgjkokehvv9U0uEIrSNnDiyvSs0u6kLAot6a5r56fUMuCOf02lBwY
ICuTs2AYOfwoPj7tnXznOS24p7YaQwAQM15kmSFJCX/czJ7A0QC51LEKGU2stFWc
lhSpiL62y5Yyv1c1KCeNIa0ZYR9RkE1uSDvIw8wC2hDyC2L/zjbfr/Mg4uOtKl16
F6gAAE1cYGN8WiqudeolZXeYyae0niLsJ5YhJeOuuF6jVV0Lbf9iB2Z8gwXJGJr0
EzM3waX1PTwODtbezoQi3CNzYQV8XZIO99sP/sV/j+IB6xmQ/vT3fpzuZMxB1hJV
OyeUcXkXOVfRyUUP11JqfnQQXnDe+Xf1WprPbgKmIYJcu/F3QwCcBZBdIO896X/z
O5j7SJu4fsskKSEFaClwelnifEoNhk3RunulX55zEiZXi7Shp+wf18hXLG4kYtUi
ybPQbbu1azgcnXPCuXzskpU9EJbcad6BsePwPmTt3g3qGhUI1G7TX6eroUJSDSi/
Oa5wDR74S3pc94pXqRWLLTiUaDOHvCR0mVaCzsWSb2whYETzoqJJhZrov++WGUd7
dtDhr0mZpCppw8ZUMBdb6pz/nvbYoYsdckDkMd6r4mlAAphb20e3HOcrUXMgKqQk
V3TbFUoY6nwzGpuSBiJ7cKlq7vb7TWxbHp3XE8ROyi8OjYO5uGTxvcl6/3E1+n1h
cNZXSbE4LnsB/kRxdyto3oB0QUdwuaB/c1HVcv8h1i/9SUEgzUEQ00CXTkX6RWWu
/k8y7B+IL2f3dhlkrOVStd7rKW57nShwczQEokrNRI0IuklSlI+JiAONfD1aSizC
5tvw7Grms7bzCx+MZ/meVV5MZPzD6lUd0paF4Qbzx5a2p8x++hP4YtdNpuVPWkbn
N1wrQW9HfV9OPVLr3+oq01iHNP6z5QDzuqt+fCHH+Kht2lcqqxxdrZoa1WgAcH0y
eBHaWvyagDKwg8BnFuoL+BTc6NcgchHE+409VBttbrsvHgVsYiMpcJgKTVlAGM6P
NXRndYKT+Ye2YyrJSy4Ft1AVjH6InFLWGI4y7kEISB1vjLxNExRS8n5y9dt/RSyK
KOK/spwnMbJQLZU0l4J8ulS1zIu5wUisEE3eVer67kcgjzuVIROBD8BxfmMOUKw1
5NEU88+naTBLMLqrEtqL11frtEqapz26+BjvNmgv82cwUuW4+ReSqfH/6HD5MTDG
xJmefAvwBWJ+iXdG49CQPYlBiyW/jvu/nYnixTvCARFy/kkaq/fbceLa5GjIS6RD
nhk62vMUCS7cGX7wRtaxoNDPcbcFfpO9jELFdpiBN4HNRUCsM8fHqtWtXtVrVyTP
4zlYaB9czMnOkZ7E3kFyTmWWZt7f71bwSEbF7Ug1FRf6D+4JDFEWYHhLr83Nw/ev
vCXocdxPuorS69pDYyLfFkJRuUrGue0ZKGWuv3KTzk7HIgCNpdARvgJ+IOYvS23K
h5gE7JYeD9fld90NpReWzLnyrbMf2f/SS2G9tsvlwh5l9A/DKhGL412gxoQH8qkA
dKHs+4rlUsHqMqxmM02pq4zVzn83v38ApH3EWKXCpXUUcZuEQ9JoSMwG9s4mrQOc
TjUDHe6Qtj1C73x88irj3C5tRSSIUsW/KDdQ3uDm0Q0kuGPC57eAqkpnQ/2a9Mue
qr9cfz5ZrE6zqqVoBdoPe7/2tnPPlXdn/9XLo/K44aeWMbQz9JvQWW6HlvhCPv13
Ig47aZZ45ONGxNHIvRFTeqAySU7VyWNQXGtmPcLgJeoldOrHrvXJ1LHJOaw3Jtu9
DbDtUrLH7QOXuRk3xBoxXOuhp1cWmLOFL2zmsplVPlq1y0MarMCVGHChESPlZZ26
N2CkEoCqnqz+tJBxnMZc9LMx7as1JL3r+xiI9/LkHWM5a/YHadewZ8SDy+byyfnf
5ufDyjbwyW65Jnv5125lm5aKRiVrmHDx3HlCAIWmtRsb7IgMNCwzgRUN+gCxhDRh
AEw2l9xC2ZOgLcDV5FAXz65Kx8rxk1XpNhZdk3PRMDuc7qc0ySoSs2/qKH7MLPfU
ftk7vXcn4gBgTglbA7LvZV8DA+sUGqvI71RTyJvkddabnk/sMj4IPY/vGUEU4nPa
/UsmTEKnrGUAiQJf0cKKlIuNBdHJW8i4veY8HbWVrlugThfEmjnq0rQMIjmuPUGv
IB+uH7SxKnugB2MT3TJkFvGpHbOU3Bg2P+Mu4jH0Tz+OgYhwuvTIcBoTcP/Yctaj
JRoP6dGrSRZZ/wreIoujF+SWiSH0SI61J0dkK3kxVSqBWpFhUeezgqTXLlhnBSX8
b7Mst1O+uRL8eEAyyN2xlbkb3NTy9iescDY7W5oSxzqhFkERfxMTa2RL8aSJ+QNJ
a06Cnx5VVRemQp+yEygX6P6bDtKt63hiA3BOHdROMg7z4MAwyxYsjGZGhK7Hk7zP
gT8qK7vG2lfGETsumHh+MEQ10nr7yC9o5rnM/K8EQFF8L2YjIgziFebNhGQmkuCG
j+CyzbXaCqcRPpIpjfEBXboacwJZfm9M4pqvKB/PhLyG47u5DpDt9/yGXvA9NhTl
DDllmrf0857A5e/8cm1tbAdR1BgPbON4BuY1BFEa/Ol7PamOm/cWkDQ34kmKJFed
XKObEFsYZ+11he85DMK55L+5O0qWIWMvt0qzBVdUYNLVVCe4FUutnhWNeUrXYO8e
UT4mzOC26sYwqrYrRjrJQ0y4V84CM00MrMnSUpYeV28asVTebsOfYz2Dl2ZYZBO1
PFXLIJBqZL14hcc2X135Xlis/F0GOceWMUH2vJTdR7gX5yU8Z9oT6fbqR+OHsb80
9dcv53mU4gILevXMnfzSEHGCPXjw2wDIzDW5Y5t4zKEsNREa1KBeh8d+Wm6zAEoM
xc+MHkRBcZNKqkWKKleXyFAyLzrTbNSfr9avJQZ/gA4WWgUz1Vp+n5dFocWGGdD9
xI/qhqeQ8bWVBUeEq6vKvo3CF2/vxrQchh5u9lhlbpyX2hS3AWtNv9FRP6MfURta
giRX3Rwj9IQnpm89kMvihOu7PTteidlrI6UHHH8tIeNxA7LYx52PxXG0p7T0Lc2F
MuVH6smakS2zrgNnym0GmZ/IyQM/V+qhalqsv7MhGOUIp0v4/beqc10//sKXuxUz
em1Wa/5YRQKuf57bM8d2n93afcAQtqeTvnJ52ra/L388aqNLPHhkzrrpmYUMHp49
GdOyA0b06pcj5T9Rz/2aOoS9d0ATMSFFk3iHJus6hcT4I60lTK6g6gkSmxCnkC3y
BfKL4+WPZINrVPobsJNga3eDLT7gKHgDGfxpaahtoHV1i9aNOGU2C4j1v2dV7nNt
8/gsHoxPW95oEuCq+S/lIN9OcH0pUl1KWzYCUiYiflbKQQ7QpH8Gyv1c6pQdrMDv
4lJQj/JHPWc6LAabLu8eKqqxLujrWQdVyIW/CRt3vp5DBg/zqKF4TFBOxO3RenlO
9cad0nx1Z0RlTk6VRPQlA2z4N6nIqDGxthrOjLPOmXP3VycsdR5/+2nLaPCqGkGm
aVw2Z+BeeZsk59X5+FIimJNCO8s6Qwyd1k46Tfr+hxAVuAXBg4GCfErCLb5Z1V0W
Zpth1d4Et416dK2BFHgaANO33x5peHUa6a8ZpNssUN7ExNhskEX4vrLtRVQEZ2kc
fu8LqDETP+fWeRAPj64j0x0+eWkiGjtaldsp0IrEeScxXFGtn0jPy1bs/jRguZGY
bclvz5IIf09fDtUfeaIOLI0a0tv/Urgxcc+kdDZ0SYdzJyRI6VZyJS7Tm/gzHupm
gKsiGH/yo/nzK4OcZ9mcfYn7FzHoZtJ/FgXUO+P2TA9zo93V2fGf8/jW6qVs0u8z
ny/MW5Veos0RNDQGFHstDOrvhNVRomSZEuAKSbvt1Ybg60LmSwQpkl6qqgxBOxAT
xEiNTX1GW64gwZDfyiXnOGSvxfUSfU/1dehCDVmKKwpQhF1NKdYgVFe3+WhfwztJ
RNBv3HLAKHuKx6+z3W9iU/7Hq8ne1d8D7g9aBlKpPRhwCcDcwG73ovAa0NxI70LO
U3UPsQuW7l8suiQPKKU/yo+fpvuCt5bbXqalFZh2t6iaebCAvYO1o0yNhP7u9nA3
JomxXqT1Ej5LyYHKr6VRacIB980QFSfxMWTresxyXTAmMzAOTtq+hTnwU7mp3R7P
1JfEY7NMMb6Q2KEnifVnPa3dxfLzJCJ/894e4nxFXbYJ5tP4FciPbmCWAy94LBUK
IU3FEJh8Xg5XozuzMtMzmK+Re2TFe17afnMn934LT6d8h+FQcnWf05+2NGCApHcU
U8Hg7W2zvsd+vHQRZOkPtqQbEes2IVsb0X/F/1hWSybpsWzh/PyweTBECr3Lf11i
B+y0yoPOdudUqCy0qga8T3cHtYo6q6vjH6N95ONv+1w/cqruDQMwLWBRxODZX0nB
atjWvtm1P+o6/BMfTwgSOIUXO85bYBjQq3Hl2VBXe0czdJSNX0chPxu7uqJVGA+q
Q0YZ8vBkraxNfvl6cdNeXxI5wQ6SbLPYJL2Ov1yXYpdiucjzUHJQPiiO2ZE4rdAh
S7V/hx0+7nwKjKFySizeIY4Y/9/z4A8Fbkbni5zGQf9Eqbsj2TVhgrT7VQALrZEZ
8Paa0i5wHEE1UVWu0ECbvzN0gXDz6+3IU/WWnoKS1tHtc8l03A+dhhw7bKkwS6ej
g7YIR+1dFQiKrAp+cHD5auNUFrM1vnZsiPwEAcXS4NDKD7XqMHGXlxbroeh1RZc/
QySC8Xl34bsaZKgZq0DX5jIFQWrQ6gRRuRq46+HMsTdfK0OW6yQ76vewd2l8lXVB
MkQRl5QLbWNmMMIPqf6o3ZoC6ZcUp97L+zoB03wPPUD1z6Is/qUappD7PcUtMTJS
/d/rP9XirvbFOQtVvTMJW4j+vY/TIBn1WEoVMSdZzDKR0eKNyVpOnOSDAfwN/j+1
F8UJJmfY2Sk0qA163rr1IHnHVh4Dis8/qz6cJtDZQFN6T0HdMicWjsyjdP6fqcVS
lZCIUgV4WJa1GGB3xtCQ64RbDl+9zF7VhKergIJ1lAOVDyBQMydoM5NzdBJ3wPmG
dA7T2cdYnm7u0toi7gERc1adi5Zt9AoVC9vrOZ+U8tz3IT+VSBMqEXIG5/fwWfBl
eOBctmMkm40s6egu+/LQ0BZOzDDSitppPf+Xb4BVMjMlnuBO9DiISeRuXCokt34F
huo08ri/oRynOaCM07a5p+e+assDQpRx7Vjlmmx2yUIrjpF2ipOMsE538pIYtvTE
tOEHNx7W8QMp/2WNjj+VgY8K5eyWrRsdDK0geUIc+wyURPOsV5sgz3PpqodLmbKD
vBTu7VqnNIkWTeYS6v+0dIKUZ3dbkcUZMUKKn+VmhjAcru4bcAwMJUoHCrBtxRBT
HWLOp8Il9QEUu21KEMsQJZM0/4kgC9qCfOJaXYIDpQUh4iZAuMC1sxnOWD4Xr7CT
lLYUjl7g84hkbN7AZ2CwyhBre20UilLQXv+filt5gFiw6QLcR8di3jQ6WSSxJRZN
g8UfgzAap6zEMXbP+HIuNjEcQBwX3dn23s5ZUBjb+Hf3Pw1onvVUIUSz+9n6YHIW
pekEvGpsnH9a2etyoI8Kz0Uyxn/Al0HRsl2p/Jk/TlXVuxlLbBU/FE3VGWBaRF5r
PvLRlXCKWw47Xse3hIdX8DIOjnT0E0Qs9hzGIfA4X+VkfWyoGqgMtxZ+HhisPBa3
wjVZWWRrvW3nGOs53vbgSX2ufzhbOO0IzGT1vsT2SnXdkS374lcC/og2xhiYYBM2
6DeadD7JI4N4K2IVVLghKHScV9+3SDRdWcHtmgtfhDf7qWWXO+x2LaDW9Lr+09pa
M0xv5hys2a+Zf1K5flAcUclXxkAzfTQ1+XKkV2xggkY7QJGBl8JmvBr/1PR9vug/
42DpfmKZf0I1lfR6KhGA+FJgQOCUXq/4uTQxII7WFIsLe+dgWMWXV3OqXGEP9a/G
ZD8KHxlh5ZiSGNnmMqYItspHJJQvwJ27LRWuRQ0Zq9f3PMJevMOOqznG0ayA818L
sgkq0o8s0sYIPSdiYZmbRFnCidDUEqHKj7mBZM+w7X9pj8pLh6ix5KmRNTbx04PH
I6v0sNB5fb+NwgWh5d+by+0WHMSr4KCiUp1CnUhE4c1RDqzbHZvO3hWZ0dXgRpdY
WAFhNaaYewwL0S06VuMkEvodCiUHWMQiNI1rsNdHYYyjTH9QvEA0NFNSNGmtMssb
7t1VuSzFVBABHru+NkmkR3JZFzynh+DzkwTLlsQ8Dn/AiCHgD1cPuPCWp+kWEVEm
LMuJjzecihvnWlAbdSNjL6NyZMKDkLVEIbdNpAuVtTOr4jdg0cUFe+eHHBXttWrf
sy4sqtNP89yoCIjvDKYzWDQkHGwY7CH4ahXG+C+SVD/Dqyv4UdCZFFjzFw7HCqSf
D+/d4XSdOYG/RuO2UBabSgeuoU67bVxiIGXhka8wUVES9+6LUOCdnCteNF/l86vV
4DulhUDMZTNBXRuIT9T8bNAfAT2RY8ws+IgPZ3pdY4fDTa+qSd1hyc7jmFdgcHYT
NcAcS7CSV2P/KLGOFLLcDBZyOWrbzPImiKZDObpEnkhvW6CaKoO5LK8w4exAg8E4
+Hgk/ssG91iklTRY8DOC/6yR3wgNUSHUOMy1DkBUa+8FT9UH0JcrJnG9PSwuXz5n
zMQP2AYhk8YyN4LunNx1IlNQsPCOw3z6LwHL2iWaOw461MRM4rWZL1wRCnnLEF5z
EhPC4oTvlIlnW60JqOSn4ipxAhNFZ06SRE42nG6t21BjrK7ZjfwBFc0JJiYk5YHS
lBshWFGeLlMOW+UIMUbnmkY2iyYiuHitkd1ZoV2Hg63qheLkzkPQIoS8qWH0Jp8i
gfcb9d+lCdBM2DOn90LuSsPJQ2/p/YUfPOlyTg/sQOY0+/JFomzWuabFxePM/KDd
n6t5M0zHU9A6A7rmBA41dEFWMKsjW/c8roDFmaEGhnWoY3Za3M7OBPLyifpWCyEL
UAUb7F4DNHho2mElD87Ksj9m8ul+j+cFN+w1Nx+2kJ2U/IW783QlIDXBivNRrUQl
Te9OZvrHL2RCR9juNac4i/eJFw0LVM/s6jWi4uvZ5XOjx0tmwxTe+AyvFjqL+GCM
ZN8mTc2VQO0pACJ4S9m8S9lYHR4kv0LnxF+xhhhDIcz4q5YaoALHy91qt8LcCUr3
FYjnbqbWKsJYv5snlR8Uz/wkyWKeE6t6w27r+tgmZPzeWqpk+KtqJHgFYdaTyXvZ
SHVj0yiyy22TK9slXIItX1YpXcqABV424FjverzUBmyW7U2UYfHi5mer0i8zT/4u
UhPqkbAadThOyQNw9nFhdwWOEqOPRnx9C92XQdqQwMofb++hYxZ3TkbvHpapad7u
sOGvpFNLEMSZVTLbopKGqfMx6l8zG6spY02UiVQ6XIogRHLAR8+beWtS7GWtVMwL
7mr2uViyiFKIA9VmYjmGK6PXUTi0WdRAvYSs/emiISR1+xrmZepL2IAWZSDsDQK/
AChDMEybbGA0y6PIqA0eGnBqpvI9qMosX9n90tiQAQz8UFeAipy9/rBV+r4mGoPL
4pGZ1Vfq3clDJAGk7DeDQ1Pt3ccBtRGoX3ByOCUkFanqrWSnSp4Va/5lmcJ9sZVq
MwtdtYcI+PJmqKSuDNDXpAnvgnqvOORNzwhTEALIQIZ1V3RXjYTd0hcRkOANVEGy
EnXnj+KmrpdWcjop1dj0hZqvCk0Za8QelZe/FFC2U6xHFaJBGgBIdgzV2jWsDG5O
NRyc/7cl8dzhJ3L7Coq8sQ9LsTkGjsYANxH0IiPKeU7qPQOTT8C5W1GxBtGg9UqS
QFSDFRIqS3eHQ3jVtJyAF2MlaB3WGw+/Aa69mNPQpqT2FQ2AUp/8GhjfOvCWie6/
mxCsKTvxuQjQyb8XfWeVz4zjCb3NVqcA74L+uMdxaia8De2EGmUNHMOfKZSiPwi8
ocpcRzp7LE8boQlFU//totoZcyREML7EKslIzq3KDOh1e+8nPspsHI9cdmU2mANt
JLDPUl/1I/jW4kzTDzvY/28F2j8T2F4ua5a/eTHIHgebs0pG3oexef1qJ4A6qXxn
UWP3w8GyEZsPo1dcw17ufNFtg1p8PTbr5ndDL1tLIJxSAGeNYu6pgXkfLHGXISQx
9ecPKrx80IhHh8i/qLXuaLqPchisPSdBTSNxq/8mxd3SpP8GolTTacYqd8047m1X
MFLf6yhmTw/E+C4hjwnR5KfF+UgqJ95pFZJyU6I/GTcLTM6Ibuh9ObhW5mRckGnG
skgdB6I3VYZQPc+OqBW9wo+vVqUYDiz8ESqGv0Y1jZsbcvDgMIdWN8t3oy5uemsN
eHwD/U2dJ4W7hrMGx1nNMj6WzuGuKaRO3Km+8w/esf+qD4fZDZ/yzd044qczPQub
z8X32mBLDjq6GHQX5+eTGFHPbDhgLdfNm5t3ABivD+mZcIMQvgAlJtQMYb/VV/zV
MElpU1CgaO4sz2yqBU9fdTrnGyzuCTfGPH3u43ylwfdyv6m72AsUunOD8Gqtvjh4
b0FOUmoCrfOgMsQDiJ2+UZtH/oqZwAZlZsTIW6ZFYx+ydA7J8kUiuD0QculxZ3aM
q6UzRE21Q/9K8AbW0j2t1qVP784SCwDA9NnMEv0UES0we3YxsxGofWM37KbgkAQq
525qWA/Z8yaBlNXb6yvJW+oSH0WMSZcvmOSZM4BdxvbsnpGrfYXtRAZVMiN/Fzd6
n6Dd9Ymky1oeUlK4mHsJH15LKA0epLfnIT4eb4SKFcpCzq2h4/gkm1lMv5mqGao2
Mml1GhTXG5NrHgW3VP+wiNwiJ8po8nMBk7ZU8j5n1EncNmdEg8lAjefaGvstEfC6
VBVCEu3pa1me1gwZ5sSdfY38ncH4Y5kj57o103+vQ7/V6bR1yjYPL3ITeG3Oa8UC
BO6o2jkuk5IPIvFSN81h5gbrjNEYNq+LMLN3WXB8trYUmOPT+92unixceTWp+I1T
WeNvgYwO2tWn++eo/FboQkYcJ8j3eKEpRe3ORRbRt0jXurVs5ugxP+dRYZzv5F20
ccLFjAOFGaw8d65J1dg0lVigevVuExJKNUBYGVk/jh4ZryMS5sZG+WniMeW/sjUP
wvd0BIwbnmHUZupqXq8+uTQ2FftWSA1Bv3quQED3wDrbLiwxaUMDa2e0yfhyxijD
qAvHS834a4O5rM5FxEXTA4RgDIdUZp9+/Y0yycUdn8eNvkFv3a7yJGIdwUt90nVs
cpHOkzcaUEMLQ+1/5fDdzsLTSCJcVmec2gguvNhRbFTCjWws8koRujqIv9AGVDZ+
1EdLxR2PidXgsrV8OdD0GH1+9MeebWvv6DWRCag5V1dsf/17PdxINh2GzLQuX3d2
iCibz9uhp2TAoqofKJ4fYkK17G4DxEsvJq/d+emY7ZwiSD7ZSVhHS1qwBdEdShuS
lLjzwTG+Cl7i8b1BDhJliSciZliscoeVWH5fWLCsxjExhK6QtJ0VogbPK6FRyXTf
7oGxyPoTOBuTqHG3kD+XL5xoK4vyVyhdxuujzPHkohWkvqOY470o0UcH+I9/V0EP
0XMIEI2VAbJ33dS8J3BVHGOzSJukVXshQRSmJY3INUAW6+6AyacLtRHUXjRbiXys
7FSSlS6zgEhY9IMVxXrWGmD9Jh/R8tBV3J6fGXKoGpcl5H1KPupZSvPgNls7xGnQ
Sj0dsw9s5Ooc4DqSHhges1/4TZimJ/oPJnKOJKmivYB7ookGyNuxPz9hu4Y6qn6V
HJgqL9+AMLVveCurNl9apk+Y3xgiRgcMxMLE3mKvVvWRK+o4px7FczbfQzuUEk5s
Q386sD4zZkXiLFyB+iLWiOJ6O1hkhQb3m5IT7RVpiQocbUWnXHCKyEqVRcoNeaby
ZSZrsOiLoKrkZgWEFWi8DtV8PUJBEm/p/Sb14hsn0s1vfCNIVztcO9O6ofhJbjhl
nmIUBNyK/pnxaR2UVOFDuxl+EuGZa05bSggDr7lvMB/VBbCfeaTGP12wPYS/52LZ
dHUx6xlCBIQX1ug6llqyocCvrIhvBx0MCdorA8GTcYR9dsArJZCsEE5amYrGbwDk
g5pmUbY8ZU70z4OmfrQiMFk+6C6+MOWeSohQNDsVmLPnjCsa8p+rnQ9N8+CV3yn0
YsjhWV5qCsEFk3sGHNXN6go0RferYBUqUbZcc5hW0F+qEG9Ne/7OlI69PmgYkG5k
vZJxBpG9ujWKGh1tsJ7O5/ESN9GHJfV3rJfk/+uMuaEFmek7TdImfhcbQqngFxlx
Q6ssF3bj+N+YELbPi+WbycxrAHfHLuzhkoNe9hxZYfhd4yukkAWR22fQ2n35tPFF
1X5TxUv3aNxrlF6uTIjheQS8fcxnPITbE6X2bCixenyeSXq/7GboSlzNFBJ8qpcV
aGWruslXskgI1XOf7XDu+EJBoRp8coE36Z8+lhfqqWq1GCu3XyZ2Oftk68PYaQf6
4AVdJtxSJ3uX+WDcVM4F65CmkGmEShRyZXjgFcPYw8ah36wW+snNh8YQKNYRFIOs
/MyZHOq7VRK/Bawc4IhDc1vnm2Uj5Tn+DuyupUzevgtbpdOauvr+qiDsV5cxfBjz
hBm8Hb7QeHvpR+ZDpNdQYoySZP/JFyyE2ZychpdGwI+dTHLVn2e/P1e8UmbJX96d
OeeBu43qydfwAjVeburVpn1aaM6RhGczUKhy1+eHRCsbp0/SUTzyCkCqTUDgTmxS
FjdC7b+hWjv7RI1fKJDyvECU8nvHiCkHGV2biSTAvGKMuBCiLvQ8lYEMvwKDta3r
hfqyqQceFm+GtaKSrjY0SGAo8I7k3MYi21CrFLUqSvLBCpoXJdpJf1ygX9tr9632
fGz2GgKN5ANPkV0GTbg4+OpzXgAj518Xn9uOe/hIyYqEO+eRuaHhA3u1j2uMSJVW
M6eKCFyBp7yzAhNKICKGBf/S144KRx8FgvDH20CrdY269+Cnrf0RC6q/hhuKcjO+
zNXg1OxUsBnzfC6b81CNVm1LUFVCeir4Zo2zNTmBBkxgYzWNZN0LHYfqWyCqKnRb
8MP6yjTnSjbFYAJxk1zmZfUkeDks+VMoHdIa0K1f9CN9jY8wMHa9xJrpbQ56FycW
cjIrKDqG3yLOZRk20JyWE9sMdRG5TVXqGnDeoMpTQ0Hl9qSrwSBm7sl4Vx2lyGxS
2ARzgGDnLUu67N0P/2mDl3TgRUFNbivk7pBobROMmDTQKZASuaOH8WhqxVdRFqdQ
Smf2aLstREJrdTANpvwTdZrnfTdr7noNi1G6AQz45VwUlQ3kMAnbA6pg7rKw6oXB
nZTvzsg7hBo6hYPa85bFEEcIgp1Wt79WJMlYv4oghOJrjK4a0/ZtH2ipaSV2Rn03
ZYGkXVaLxejauVFNLPz+Ajh66Zf3C0vkjLukwnTXfEPqKedWaQJ3LQfGG80qFFCN
o66kfp0H4vi6vxmByRIeAYh/J9VMfXe9zaSjcH8Ki/mfMdPWF0WSHTc0Sx5zKZw0
vjjs9CwMrFlKA1pRIkPqtMi34ZzalTtenkYqzat3TMyFcrVsnmm5aBf9DUEm8rIS
A3TDDRcVIvLfO9yJ4XakKhqEcbK/nz+u/Qk1aIYpJrWA0rhwFeJZ4iVgl2hC8zuB
+gDkUij9iwd/QBLFr7e3+8z9z2zlUVk2skzCcrgyaQz34rXb1VA3x2WiMrNLWGpL
RKPe9ny9Yw6QvhVk0h+P1qfX6g4DOixQDOjSMiyYKqa7F9LStfiHR23oKqKXyATO
qCj+F/SHRBbVcfbSXO6fdSG2urziP4nV3jPp+KjL9BR3yhEIvhJ8W13QNDeepV0L
V4t7QbLJ8Ort1xyE4a6tl5rUdDuvT5vx1iWTDzm5qu22ltsEqCLSJDEltZOg99Q6
fcL63rygTXvN6sywooUU997dti81AdtjzqFqsIxyfbfQzwYMguaM5KeW9R7D1a/d
zfVLc/k/UFXrO+fRo+kzHYHPIIENUE2CY+eMUhIApe47cOqm9FsGP5g6ImfN4mmk
V4SsWRuTNtejAZssreTT5fp0hfQzUQW5gFcG0+mbKe1LZh0huz/dxNIr13ETGHkl
TehJW9LUjATkQ6WGc9juNA2qC/SBxsbtlL4Tw0eM8a9YScIE4gvnDrZLJGsqjv8a
8W5kYDwPLv87OcnrxXARbhorWpR66pV9q2Jc2dgaDdBWAwGjXwbFwjbQmMMQYryd
jyzjjWytW6z1WzNmUFuEjC+ZhvWY0MTmr8xfypESZgLATHTxd3eNKyA1lRoJ4EdW
5NzF41/NNhVI3gKwnKZLn0Zev3lEhGzKnQ6zYiCCLRccLjMtWHbAoCOFAWMb+IYw
Uip0XBRdjtgzxbXFIxSmce9LTe+iunrIesvHVZH64GYtppGPd+pUJ0noGtQut1u5
MP15fFzzIVdEUiMLMnn3TO1YHAr6ZOnITzc5zivJdx+SuSBKAPsQUQPh8wePjJr0
smso1erKUgXPFWsw8wr5nMXJrSGguWer2gcSMj29QRH0la3uryNgeG1LLufYgqn3
F/U+Y8tEuZXQJcjzbSoQ5V7IWT5iv3CWhMb53ZDgEafJkLzfrpP/BeJTrZzP+mOV
hl+l1ynUofp5An4G5Pp0XWUATv0ouhLSEfZn0eDpPDNqRKjm+XcJxiJJTbV9hnQw
+3oF6AZ7q4IvHxVzse1AxgGqJ5FidCwdH50LV+0SllRALtnOaGWGzux+KOD4NfKO
pT2HIlaw+ZzQnUQJbQ2Ue+665YDMaPwJ4zK8O5+ttY+cXSWkJ3+uxqY6p6s1y9Gu
8u1o/BDWmaWYX3i3vsjx/e5gSt5Gdam9caGUT+w8v+oaBnSh6Q6Ps9QJhViY+D6u
DnBtDQgIc0xsI1yylKqwJCej1/zFOW+hciNAR5HdisbEP4+OkF4EKRYD+jJT5/CZ
x9gDBXcbPf6iSwHUUkTr2rJpU1U5VJyRvtq8n6M7Th7vi/HwCYUVNAb7RchUMOeR
NXx6GTv81S/cgbA4eiWHi5QdA2wAhrhZEdliqMKipbBEaNNhTpnMiTMfFtgfkZcT
Udqck3P/egmGwO5Mfb9c7Xh6mG2zzQ3yWoealvWeqUwA5mbv6GiyxNCq6gu7E99o
vRR6otHo/6pFgI9Qb/8m3XdkcZf+DGjUB6S5XLxBco6rR3oxWJmG+uuO6T8+U28n
FzIqkkq6mrjpCLrl9Nzusj8U3pdppgnAI94orDp/3P+hMzP3UwgFupMT2bZqOj5m
dpG4fBXpWwULaNnGDxbxriMcmMnIBCm8FRIGrYC0gvogP5JFz9eF+5F0WUAxyBog
+lu+nJVhHPwYBT7SI2rG/nWw17ZS4RP/UWwPySLoQwRtVZOItNzSXMcyEHEOYxen
PNHacRiFwAfyYri/UTapfTZZyse+WYsOy8jVgpgDm18LIbefhmlW4EUkGErJpW/t
v/LySnxO6vu/QF5xEmTRMxk/MM4FuGPcBqR7NwvDcjzApp60Ji8dUExmQqwVeafO
664BCm9RU/xV0vqgCGGG8XEMi1DXgiv/OMeZz8tZ801CSm2MOzRoNm0PsHlncsbN
JbtfHDyWj3PwmKX1b1Ru9u7cGCQ7etZAe0Xzl4lkYI1BGjhH3GNrAi6+onNk7ajG
Ggyr0iyrYJ7Kw4TDIpL7lFJGBG1ubginaG9Eob6E4oFw7PZjtaLMpOuta8iWOXTd
Ktrrc7WFKrp0tvZ06aNAJ8wH50qOebylH/zXipEwKq9FEDd+4Yxm9ZnTeCywfIUb
pHYNIoO8WUnxDtl4SlYT6Bkf9Gkui6ptlNg72/OI/dGgGvgk5wzMHE3SYD12DWI9
3Lf4KuMnICMIesRYBjkQSFl2WoULozjMUkor05OrcOqVoTlq2WGwGpdRX0AFLOHv
cP/PLcnJVdS5xMNYa7rtUFRM+9GpB6Sfe43oshXfG32o6RR1fKwIKg3fOgdbZGdW
JcW8DGik2eeBD6vb5ekMYnQgvAGNQ+jzHOE7trGgGqv7Um1o9IoGAiVlPSdgHkqH
yahY7RzzQQfhcwyjcEVu2RRdq3iCUG4JWzMZwsxe7AzI/K8ZNpwpxZ1qvausqvtA
KTQvlCwsGOmpuI4VFcLg0jZ20PLRUP+zYLdBCwgnRB02YFNc180+gjqi7yoQxN4I
HKfZI3UiQDPC8/vqq13wYfNFTXeMfjZHScEpJ/20B6qzmYQVAmNJUoSnvck9SUTf
ZbbDUJPTR58eneDmxOQnRccdOWstwoWnjZeiOMTnURI+HtbWXZw8IVkh/gHKoDs3
dSsqnJr7RlqOOGd8+oBZT7PHfoNUcsU0Dj3WufG3T9AoDkUEAmZ1P/hs0lRch9Vz
5dRTmHNH6EM6y7d0TbEn52nBLNjl/JGje4rToSM0OIX9DinWHqHxGSd/umGKMWXE
w/1GrYDppIPwy1HrYkt7/+10F/ZcVaY+qrTlpQrrJitZR8bwxzCp6WiB0L8urrV0
HMXzaUgG1L4S3Jgtrf9mjeOjiPkRfGOPur6N2m/1RbMGAL7qTW/jJvAY/7pjiMzW
FrKW/hhIf3dWQWAXpWpXbGtLHT+4xdcQfsq3yttmfzFW73bnUN0zD34PZhXEhbh8
emwm7abM4avH4cG+E6IPk6sWFQqnsW6MsdgpNyPPyAVRDM+8Yrcsa0kpS2lJXjC2
ZG7THwegTHjJnBlA+ao23TPEPrLLR4eQl/D+0n5oRAG5i98Z3sdcYD0YTrLvh6TA
OwF7nKoO/cmG3nxpIwKj/ZBONjxw9H3cZqLjKvp+/0bibA44PXYsNbUhJ5xjj/eG
fiT1kHXxqDKuVvyYqBwG+9ZHagzDFP7DA77ZyFC75hCo/BAhso4SILFaedePlMXd
jSN06gj7BS9abyVG847PpARvdaUZiIJ03I2JTeOb07gAix0NK//J2ZWzr6qUZ5d2
YwmarfpeaIdBm5dlF+73mhOkEqqqq9RnGGVZH9TNsq4K9ih8emxvf9CxPJRu4y7J
VpVSWnALoLx5v0N6RPKOe+ZLfjJ4WgvQZs2IYsgOh8+gKT7UVNGyMrkhzL6pOX81
LZ9ssMiAQcw1z6S+YOo+okGnjizbs44HbIxWoisfGaER3c+s3XD8vRxVSgxMjFpe
OIhB0vwvS+J8OGcfbZ5wygbFAMyEgrfUe7IKxZyeHkLh8gRflM2ih57WLGw5AAG5
er2DVfhzbBdpTbi+WK0rgK52W93pR2hDRcQz/wjq5ShmgTwedg4BrsnuL430g6kr
pHwvTB8/5kExJeGoGRaIH6fcc4bSP83S/978LEr/uxbpM0wiOApHMVHWVI6OECGK
QNF+XrUS3Kl/Dlai1hG1Eqc+LN7jaTvQDx9VY+g2Lj7FUnhVcKLtX8vCZBnF+HEU
ZuMzhP5f9hs/gSQTBSJlPeYygOxm6quKrLkKvvky9L+pHF4QEViVcdutHmKb5vcs
YgpS5ZFBnjl19HfHJJA5YHTTdlKV9wWub173Ezxk35UEgFJQ9OJ9PvmFSsouuu0Y
ox+0PXI72S0VejKhOhy5NQLh1A0c15lwdYidKlh1uA4UnHmsmpS5IwzmvvUQXSli
D3CFq1mXgW4PqWJv8avIoubpA9VEjOqZAIT7OXNx6wtCsLXF9/yuanZ2SaOnDqxu
JaISwyYizrMy8Aj7WDQs0C+w6Mupe8GXMxXdiXyqqeE5NxEHeDcCOOxpnq5Oia6U
DojrMoGupYFgobZ7LuYDwnVx8Dmfi9ew9khTrYliY03O5QnmECL4CK3/rg06zGjO
fq3w0z7zA9ipYD7I9UkYhBmghU1X3LcCCjZMha/vqnhNd3r4K4NgV4AgUn0ULAgu
IdqChshg5qzBshvr6eRtiwRJoex2SMDXnuVT296oiQ5jHLVnHpBi7hUTHqy7AcTH
rovvRpzI4UlQz1L6DAI/jSkMr2ZNIljJSzutFKz363HiSbbNlkZoIHT8IcJr7sQr
XuDxpg1bVg3LX0uKUP7LtsEunW4gY5tRcgd0DNDb9DZlTqxNNXI8i7LGg8UUUce2
ma7EDPffsPngJkzG7wOT5zQGn+TbAy8AAQeQpL05Va2cqEXNer+tBuCxkR3eNm1B
GvQL+5pgHtp1oHNAq3LbBAazDKYoWTzZ4n/QilmyYBoOtsJLkfw74uwvqecWKsLN
esFbMbE9uXallt5osy5DENlOSksCBIcjlGOas4wO5yOBFy2ohDrYCJHkee8f9ByW
divtuzXQ8Ao+hg/ToVrLFdZtnHBp7UqSd/C5WEiPKS40QN0ZnkSRYqZTeBQq6PqJ
CuwdwumQyNEyn3/FqgX3mrBAYHoR37Sjk43rQp2ahenweEUtYGJyJbFOUglCPnLo
gFKeZyiesSktzEE1b+kNOxjrBdYGLR6brjSbblSKjVQTIN/RvTzHXupsDMWSzPiV
MTSzwa527OXKmNc++U1B1RSzM11MY2Y72PAxtVBRvKJJWQCihsCUE3uJ64ZdrB/l
UWRnM5dRoPCzcLPSmdtiYhBoCvG0oQDtnjwqKUHErHI9GBLm2gk4x3grs0gBAoOU
fkQ77JDI6a0AV1dwS0rPytO8opB6YjhMwVnAvvtWBdYwYz8YG6lNpxD7IyrnLRy9
vHEm+IBLA3V3uNAGK9DVe2Gv2KvOI3ngKvDSYQlevG+PQP53JtYtHCy1Q7RXwvGv
tbSVlURX+7LpWlAHTIrsmG5lb3zoo04TnaSxEeBOX2E0oktA+WO+Qq8EHP3dSI2V
a4ZXB7U+b5BFaAD8payFLMhPAnXQtK52hfEGjgD5UB1N58NMjZq8zkhQFbkcgOPt
DKXyPmlXTIJ3TmhAODjUl9LubMu0Zfb0Y+EI8v2I+UUZJQnd2GFZZhXOzlzwVE80
dhNveQSo0dydnQCrG/FjyuQhMXqolL6hNM28mQ9Kym/7bavVvJjosw3bg/q1eHiL
y80T0CMqWmH9B1t99DvkxlVocDOLy/w89LvTeEEGSDL6izQh1d5j2ezXUu3w+JzW
hhSOzQ0w6LipfPlW9j50cejhPEZWov2vA9XX6WG+4HqbTQkrvFp1T82oMD94tIkd
vLHUu1MUhKcDFVuU9wpsI529uzTX8iHD53V7rY9ffo4AcFtuTIIeDmrnGzglMjzX
772WEzlxLR4Sf4Gh3/8UkOcwRuu55bAMcnV7RiDTmFL+lmnz5tSO+c8M30TOHrrJ
AmthykdFuh9QXYhO2BNGhJmd0YdAXexk/mnKfx7S986/+UW9DOGpmhjXpFjnrSdA
FPuCjLisB0op3PY3EOv3LWr+bgswghkSkB3zIxdRrdK/V1hIr1UdXu1Fr2IYxB64
8qU5MEEIBKodLVlu4kIyPQ7HJvurv/8MohiDoRh5E608yJD9uMXbCiGetHWo8byE
TjB5kF0hdufiQLoIwBtcJa/LV82ZVguGLgMkq4zB+XXNl3BmsLXdLEStiFuFsidP
WESkfmXpQTdouvbC3etisGa0cyV2P88DLsZYu1fwTNA8WY00lNfxWXCscbnlwmgv
ii2nZlEjoFQO8sELikhJenJFq8mNonfPDnWctb85GpcAISJfZcywCSD4AU/T3XKT
lXFydXpLTYoBQuWrYurmkKjveQnqYp6F8/3tp8MKcBBe1huArzj/GHalIYXEsjIB
VOGxqiAwx66joudlh5r62mFLlR+Zvf2NzQpshBxbATgKySrjOdZDJ5zr1QNMeReL
ycvS6kz8bK2mh950mOEmHx3DgNTE426KDnurqFXvsnviPeXtnM1UedNTLIjnvLg4
qVN03aKuKjBbmP9NG10R2PteaSRpz09Juk2+FGAAo6QgUv05/si2oegJw2hAiehP
tCYPky0ANDNno53Fcp0eeSpBVFAnnjaXFuJURtVq+g780XtB295MbHMZTiK3L10K
PKm4K1gMMAkxvhCIW64JODzm1qQ1xYSPADHBsP4wpsuRwUHGyFL0c1Z8IXdgBCsB
cbIpRcSSugIHm2mqY2qYRqnSBTS5Tp3A6StS22keRqeYyDIlH4RirpqKeSCubeJS
9si0l1Y2tMKYduHEAvJlQL0J6zWHsk2gwnOIovwoS839riKhDtnLi4h8+K0ZNrS7
NAvsIjo8dZzgyl5rxql+wF78Tl/Q+DZYchIk9nFoEe6xh/ZVS91I4SKZQe7EU2JK
Sxvk7YZsPztWyJ64gvofy+N81QqM0HxLtYsXA/p5M0m+GAB5PJKyDvdjIVo95nr8
PfH20oXGg+RAszdBrh9KRbF9Ojz0Nq+td59jv01xn0xnlgrtfsDJSYyzovjdVUN9
2+KEv8V4wj23D/fnFlIj7T13AbC4KDkaDkDVgljNu/B6LHXyLIgR8SKNmCgcKZx5
pCkFlXg9pkaqGeKL46yH5eDyPWn+phB8gKKKTl5758tHY4iDV9vbPLkgwYUi54m2
qfATwufxzRsvg5kBEMVyTfAEA4jbYDyaZMf22veRY7zZM9t79Li28yJR4tKPPMem
yW96wXkzSmPzNVWnTlYuwPWYLKatbp++S8zWWc7Zqou1Df44fDANX25C9pLURezJ
basMj/TgvBXI9lwOeoSF1qLJRkkkhsMVhAsUTySfLwogt1+Kd05ozlRaAxd2ZhEx
1InLRh597r2Kwfh+/PzwHCBYp+pEFVy9ZahZ0w9pD6MiOcB9bHlUMX/uiPlTx1mA
lOXqTP+vpKqdOvpVfvVpihx8XmgmE50FWevXBN75704PDXDkrqfFZeGuvnou+YyV
e55I5ChGazfYkHxdtZokIGDZoQ1IKZfN1q+OY575SWStZOsRcCrCtl2zxmuwkeY3
h4RpiFvN2umCd4s9Kd7nWm8xoudmEC0oZDY6XVtigfJkX/CbCjLOrsaeI5jz8wTg
pgzaOmE7WXgvNfkNzKLzLv0wXE+4tyGCXJqIQC4kHGs6A8fHtLOtQXbyLFVpqOX2
sPIYaaHBopBNfyLtIm57DHFoJ4S7xYCUL60KrZpBe2Kudibg9fxGzX0pb/do2dUm
+lS0odJV7fkbc/C0yv3ZevHqyY8HUfys3O4HaKqtZobpOM9SWdqKN4JPHgsq17oK
f6UM+l+zkc81wc8n2WN0yKW4c41lrhrrduHFDTh67y2mrhbhzBSGLGFedQtDOXVI
pfmxKhj7nPp3MjhZ96SgKcSe7dX5QRjshsxUSMNpZvAzOPhUXrSgUArrbewQYZ8r
g9WFiQqzpA7lAvV0sch9RLxkt6ZkN+0fkpsERaPP8N91C4xApt9tDg3LGY+voAaS
AgybnXH5uf2XxAGQg7dMKqCAgAkRzIsvBRbSKq4EbmOnTlEJEqoWxr+HPmLufzhn
8cDn988tz/66mIetIcJ5FQuRw8HmAryX4gXRtigvu/pgELSeM+xBJ+as/ialHwfP
hNkz3t0rB3anOeRG0IhB6+GCBoFnsqxRZXZVN3RmcQaqTcK3bbBfbm+LRMby/KyH
p+eb8tuY6TvuFC/U2Qz+OgbX0hSqGYVm3/MEcQSdVuG7b7d9Nyj4n5PyEeApFUmk
efD9CXasGEUx6F8ear5AV1E1Aa3zaAcSmMYSLegBkNT0r3sT57wP0gBAucBj4pa3
xLebiNPrt75aUnmajuWnN9joYxLCV02kgi24O1wslRThNDMNM9Ayg1Dz3pHVyq9r
OlIJlG6eBbunjGmNcM8E7+bUqQsYvPzBEVPxGP/0feZ8W1XSGXNjTyqSGvYqA/8K
bV5CaABFy0UeKaihHY7EZNvzFcdyCjcKCaO7Q02r2M7w6cImEwlsj4QnwiYQZKXd
dUpS66c0LDVHsX7cRSa6l9qaVcsu5lMjStRNdDYOBLdIMQdQdlHA/3hKuPsPayae
iX3CQ/t+eBBQhN2dB9WhOoNqnr3Tu8lJK+p+x9myjhO5b3+2SBeu/dDM8eBpaRuj
INKx6nD18abGosn6DuMmSUONmT8aCCLm+oHsrsHK7Gdk0/hydMXGquaQOATNAGW6
INtCwsSgw6oG6XMl/YAuJBGIpAT9HDoFsv0oUteMZJexiK8UbEu70oWb/UnjU3H8
ezBOB/4ao9k/mN9M6iQctKIQjGkiVqe0yKT7i7IEc/vTT2E9ANt3ejTyYlen4sWD
OkTpTfVSjKsCZlyZY24WX0cxcAmBQgWWJqNMWIygQKM4ddcNhKrGK5DNtm6LMVRz
k4+IWN9DFKnj5EI8Na3gF17m29T4+AOjZoxx0Ofij4ggl6hUXtf7Ft24nDIXktgE
1OpXQM6bdYIYzNjg8CEOtvoOfqH0WcG5Nb/SL55/ennjz6aNJO1eVZZ7Lip/ZgQd
K3KNYIHbZC35z8WCUg7BrPIbtE5sOfHYZI/vdjqhRAF8Ftz5eKrO3SbFsWGCtZXo
+WtLrR6K/zybIYU9fOhtdHj2Ylmkrgha0r+9tcy324/K7j0LShfcM6M8fOhgZr2N
XdF5EwT6+kS7IEurR/gpfM0voURje1Tp3bkaalTwlhStdKQQEARU3a5ASYY+aNpl
5RHTuE1Rxa94icIqFjaDZQJAkpvLYC8N6iq4hykyJ6Yjw6eetCcvL3tru0vNqfnG
spZaScgfOwnKS0Gt9Kt4U/Aig3q0qXibgloo0Njyo+q6eShGX+OT8jlFufG6LcGr
Sg/BUTE6gBDGPjPivd0H89fw7vs7pRjHfsFZ6OIBI+bz/JV+y4rVP/+eK8l8ZVjg
FGfs6Op0oiLfenpwq0liw1XGmGjdQCuSV38OGQSANGvlUM+Np78qREG/l/tzJ8Z9
wg0Az3XgG1HD2vBsmB28usrrNjyVqIITyGwMWERkE6avYqesPdYs8fh6KO/cR363
DWBkKN5B9MaDCwAqmsGodEU3We+YIvEiqUmdsklR6FI5ST73rFVfraI5jOGKRmWW
KcIDlMvKwyW5kLsgfV4SA7nhanJgv28VgqeXJRMsSzgaTe0V52uB43fiHH4xEQpb
4Zm/JiAc0iikBye/FZah6NKA+XPtOI/Ntu3Y/t7XLHN+Syi8FGX7TdkDn/ANpitM
G6Bz3v73Bn0UbOAv5mInI+K0lxcVR0OjFQiaIqtc8CPLw+ABH1zmOS2W76QB9o6d
qu5SjtFJmQbH9Z1e2RNnMpHXrFYu5Owlf5BQy8CsGxjxVbnL1rBD3Kte+zylFOz4
+wjz24OYxJA2/NOOsto4mMZ/lGvq4t3m69+zSBrWfZgIGJ7wB0vDU/Dh9w9ELAFs
0J9OvfiScY4UjK46SXRfPFkapIexBDbzsUQ8EKDMy1AcUelLioKuapPjOfrHysAF
Lr08eIJNvwJ4X4YBZW51hrBEC+jYWiZat9QpSZJd5zi1A+gw/f4IgNvNHm3Yns+k
mSZxwnYEtXJQxDZZpZEIhkep8QNWour3kpyExJtygr+G7jGH9jBpl5s0hxE8VfzZ
5G8SZEEJXjVx8ZGU33Akm9Lu3HIqzstT0xC4O3A1ekIG23rCjbNz7uaaGHXbJzgX
//AssRcfqaIoTsbNeqnsxSSkmFGr+RCe7yanAVYsGpWZrGiQp8JryytE6DywmQ1t
YtvvcdxKf7SJRCoGRakOWyGqUemInPv4gmLGLXF++sJUz8Sa90/l8C+Ikp90Ugwl
Jf5k0kvmWfLWj9WLDyDqBZtSC5nVh8VihDQIhb8zub3raalhHGoRZZM8LL6UfBUJ
em68wtjy8o7HcCzCZMas6WmyLrQZq4Yx53OjlZ1IwIQBC5WK2zXLSgs+Xlf2LDHo
owD2danzKpoP/hARsfy6CZoaH3/2UdCuvm9ve9MNgX4+L03VbLiLr/vtxW/iyQ2+
Ic29k9uOH/JdIq4X/SqXPkhXRg5dw5BWduqvbmzOQkLBv/L651fWmz2QYZtr0439
ftz7Mmcygbs1UAHeUNzmdPfYXWUqklWVxJCoWidgVH8LN+sGmSStcB2ZGv5pXiAE
1WcD+f5CxGu68h03dK01rLfaJliQkzxviOPR2EFNKsyePIK2yMNOhIgEh77VD3Xe
f2O83YCU/LMCeqd2boG1cgu9w00iUywJxQ8DiDG6FLYsPodF4gjK+geXJXWL5yCM
Gpkqhqy9oh55r/RPYmStCKFYmam6KNx/yJNPBlHjlBjt8ZslDkEQO2y8JYBKGjRM
bLIWBZcbog1ivs/kmlb3V0+TkK3LWjhpb7R42Xnu2SAvt4HRpngEdPzLpL2Gw3w0
Pj4uj+9Suv9VSrxiBtrPAHgBI6k2ZAk36IwwxFVvcCiSc8LYgjudxa8840OfHqjp
17YNl8skC5xQ/2pqP7aZE8zQpBwDH4YpyVC3Ikgr4f2wAk9jBxDYorDiLdBFWowh
OputLV16/6LxypBWkTcExY8bn0FPMrMH2ZfTIUnJgaJ6Dg4371kekBmHP27ygFWY
c1Ibc4AC8ufv2DwgSuodDBzKMwcnI88YU3cgI4o+b3O2U8lskxCsGj8i0nVvl2CC
9xR1g8BbGOsY3RVrFWVLr3EPi+e1/9VaFIUxfJA6ntzPfrKXkY7dSn2WZJhwzhiR
DLSy/hE+b/SI5E7qkNpHEK4GxbFqQkrPAaMd4LjyyelV2HzuXxRIVuuXi2ThgJlC
BjOezWqf1CTtcIhes7JjL1txhHIcRPsD1l1aumfCIr56J+telntnUs3FrecoK3NI
uP4wbHksYDX47teKjV2tzpAqZ0TOdGi5VeEy+unLyX01sNTpE9kWlfLwdMoLVX7o
C6wJj0qc9gYJgG+QJ1AvMQlta1i9tTOhKUJkNt4rd+YaKuin6zmREU7T+BX7htPi
kzEA05pyVg3VJW6E85N+z5jhDEXueIkhBL99QS3MGCZ4fYdEpXvmWvwb8gFHnaL7
6k6K5dsO28+LEwHis4xCu7JOKCwwKkINChlBTmzSDeGTcMoCJ8KhMCPN3c7gBAsH
FX3HQZjgpSTwM5V6bkTyAC/hMYh+gHWkLlJWjrkthjJA0FlMEQTwCZuGoHpUi1yw
jzJAptHWmjhUA+aBhw28RxTsElg2huGRRMuNaZRdz7K/Pp7g4S6OwQhjdQFVsJ+T
xqAQVEblXqMdPCua7QhQR7O/7Mb+HTzeUvY5Elx6So+hynOq6QytbyGbonn9n2Lk
en3fdN52aaXtJl6d9oIALWfwVsPOzet9cRSmddEJmij2M2zda99j2ipImb7CZNxZ
l3SfKqeGZyRjHrthH5EuuUR26dJwbNV1R9uQt1mlxfTBQanCxSRTpApKy7b6XMFz
v8vjuOXDDBMcbJcGVccyU2VAWblOrjItEHn3wBbmfQyhaUUOZlzVtc+Mf2oSigJi
CSNglqFI4vHsPq/nJHiTVzMWISdJ1FHaFWxpjCTnIk7wwz48lHqPiBMW4H03g3Ew
+ssc0WqxxE3DIUNmUp4H6/DMRjHPn72NmjYhHAKH5zxagOmPZxpxqR3oCkGeWJEx
6qP53a4gOMv2BVCLtuiEE+3Y9GmZgAG/a5k8YIlc6yU5pTtBfo62dPOrCm1CqcjZ
oRN5OFKnUgZN27EctjpQpLJGg1zkGnuT3ZouEkX8BZdSADbQqW+UAM0woHfflce4
F9aMp/ElRgzSBDqPEW44JtVdwrfKL07WO5LzswSAGuhNPJxlvlA0TjUQ4EfDJl9i
ZFqDqku5OhJ0DUhkpAd3npLXgWSWDH1cVNMQcV7hdb2ppOWxAeS/HEYvX+ggWld4
QwnT5YjZo2PjmHmKtQ2bEnkmD6dBbc42TQIPHbTfrJxzISRIwvJFdtN7W2OII7YX
qWIVaPnW9W1vd48qS3iAVQxZNywPn4FXkEoixkpcvGA6J+aW5GTgpfQSUQVbmGag
dFlMz/6wKsmvCaEpjZFAV/MbVpdc2nDTsBRAE062PewnsE2XPj9PByH7Nc9cAt8/
RJE0KANWdjTnNeLm2Nno+9KdWDGfWgOBJUWhyFveL5PBYBIIgd7ODzb1HEjT4pnD
/fkPakdyPLj1F0n3qN9CsHwiMkA+V9/OBuD6KYd8ejC0TY4Ndb05yGeJQcKF9DMK
OAiE26Hz2e54LFlaMKIu86ZYemH78VTEfiY71g2/nyRHi295511aQwdgaqFALPaa
f7WzeZml+uZ8AmM3hG0c19k/YM256Ap5a26tW9Ej6tcXWSAqaOhUk6kAxKJ1v6hu
FVjraMq3j6qm+swnBoSkgAQkqm5hqOWb7LNLx5cqO7Jq35TCTed5yo40ZeFsV74L
FLfiCtxQaBv9gqX1KdXXvFjXtZDFr907YSdCqG/1uz7Png8PuHWt5z99bJUSLlDB
zQ6PMIQk5sQl/N624Y06ytIUzTrLeHpwr6jVQNx0D+PQxGk7UVemDJZtyMG3wcSX
DWjlmc0CRecWxhuvNkZVCDo5LLcboRUrrBoHZnD9tmkkVbTG6+PZV/Ov3wQ9CS0T
S+Ha7BLRvL3ptgcf2X93tZ5kf1SRoDS3kTk054Isc3ANM8BUxxHG5EJABx7eDxAE
VQIfysp3kHG3r5umxd9KSK13M0yNbYaXDn7twXvhVqRJDE64+Jdu2aOi2NWeCRj/
pSxWVrtz/yw1MQ5kkUApslXAHQWVBTgheUrc7d+GJ65VCsm2+RETH095VXkI6t9U
SepOY9alLeBgmsRKhkr3xk5awdvykLbmUUrSSW/HKRP/jw1zMStEHWBbGhsKBezY
I09gfM4NDFKBJqANLbci0CAxE6poz4VmUDBdBIfpA0/Umh0VpCJ2pwf6kTQu6FSQ
q0+VdYrcagBdRfZLvYKG6eH2mcySy8soXeYMwDnO9iqnHkZOFcQx0XUWkXbirX0Y
jp/Yir/7Ri9dNSCCE3OrIYPABT5N0amwmk9o7mwbGtcbRPDKrhbbWDRcn98Ro+lw
OIFAZuC5hWFTm019faRwfAeEyOx6CMYuKNSjcRRX7SsfVjj03WYvkOvJ9xEVdRcs
t4U9UI8urPboJuZnE77rn+X+DDGxi35f+/WyCWfP7EocSzQMy6QGzlag7yOvB7YI
CLxDBfleTmoGhIKkJHejtJ3N+v8mSiJdNBnV9IZh7rG7GP3j1czERhTpsd+sb4cS
QcjMaWlKmvKpDRQquKvK3QebIFfeszzbKUizwKAIhQvkEVEgxWz3378ah2uJcJTQ
V+RhZkjMUgRYVy0/H6eMvsyfdABfFqnxlnLNafD01sX2MqDfy1UDswdl8XhwZOfb
yYDDLhOW58Z7VxVfJJes5vfDQDWqUm/tPH74LqU7lfzXHXC0w3WTgey3PebfkF3v
zttULyjAwjezlLZY0Kuwb28ccMhSX7d4jrDK1PPPTHp7b/WoBpOvRob7QHx6wudn
zjZJ5Me4r2LtI+jf4g+XNYjMfbz3HzQVSgL49Fc2mitgwzew+JxBFXhoLmDYd3pp
HNkA8rTZf5KExcaf3nFY2B/XfN2OqPpNhH0W38wmOZiiZqwXZkRMhTVT0G4oI5bE
9C3OoxskMYQENaM9iyyBuBzyXk8jP5gDFP9ByIGN3tZ9qqkjpjNPUn/znoQUcjzQ
fVO0YtYLYToFkkwNbpHb3P1sj9ZQ/aCZ2wd3wedHI5KksVe1oTlJLGU0OZz1x1FB
qIRrxFEgD5xZlsYUk8Jjk39D/kBPkHd4s7j5CWDWNMHNzVZxiLIk0iY3EM/im+lU
TzeOSyejUCcyCeu0Z3zJzaHLd9W+MofJyPqS1JZiYtxh1ZuSwyAml4Jk1uXtZeH0
pLmvsc8FK1NNvQa2mwwqH9qI/qlgwrGzoeqZ/hpaf2qOO4syZOCXYzYQn8U5eKFj
a9Bx+BXPbjqa+cmw7AtHnUNWuXUa21mH9XyLwZORo7Or2G7R4Mf/iL+M+O3MYN9t
eo/rTy/QRW0dZy5HMV+lW9DBIurc24NDsYEZbSqMMCOPxpsNviuNdgkVNO+5xIRc
r54fbs7NgsNjlEln7671lPFkna8Hbq6pIeDVL27yfIRk7ElSHt+/wWZp/enW8567
bo55yv+RPQMQsKK77yUzmCgW7HLkxaOLo6J91kN5fTFA8G3gsgLzEH8auFKBcQjg
3ZPTVDFfxrmbUBejbBFOZvnmMycrHlrgV0CKnaIyXT9HkZ8BbKsyIyfq9uUzk1Vr
TV6snJ+uTXWpFXXKZAdGKmSJrh5BAxggVF3UmNvtQzQOTwGt5b2xompsPDi2u0CX
6GgzQOvtbvt0Kyn7qUCMjJrRYqJAIizy0EGsO9YSp2CBNz5Mt/c4/HndxjX5wfCf
z9DDcBev0KQWajo0LtkTG7yeSbMVNSU3jnvsGyMsI6nfdfux3I3YO0itnJFMrq8Y
4V5anky4rO2QmmiA0mLDEm5OTbLXQdclnE22geqgTds/hjguu8L7hmAzHCFEAzqe
TVrzYWirguTT280BU42Xm4KnnT4gMl9+t4BcEfEH32sjdBl11dWXeOqi1kTycBwp
/d7aHPx99r9FXW0CNQKrTNlDZj5k5vF88QF0wQ5Cd2cw3/Zum7AL/8V1xheoK1S0
kfBeDXbKocV9OjLfu4Uq31BhkzLuD1DPcb3MchdMz8rOWOkxKvFzcKX4weP3FyJv
s65JUEwQyrzkZNh7pV6+y3oEn7dIFkf1DeowRmXQN1Y8CE3H7OctJ6jKZeQqRDsR
tbg8i/BM1nQRXvCYakZsctyb8bz8nxkRB+8DOs745hG/rEcPQ9A+Q+wbGerRF13h
yi/FPu69kLXUyuaW57ecgrRLAfcSj9qVGoOmkNuJIn+TkXQH1KAvrMttrFk/CL1B
GG03M3K0NsqBmJOuD1iVF7IUihWMD7LJetGRyqL65ISBnXUuBAQYV+tV4S5GQjco
nuWB7Hz1U+se76z3Vak+M0YlNNwnLmu7faFKSIg4wRHdu5hxLsSv4QXiI7OaQwD4
HWTv/dpNmQ+0tLUzeyVBMC14B4+7cCfPjY9ld100AL8uVNSbOfsFSewqBaY21AUp
ywo72r/K9uII6X/uX/54mDEhFJFpWAIvjYxdttHRGJrZbJ9Tjs8DeijEUuHis7BC
r0CRJX60s0eLqjUOgxOX1gZxWv5MBX8HezQjbCThmYlmxHAZUDgHA3zIid/NXEvh
VbMFpiKNW6SjV4JOwii61mO11NjB7Yp1HReI4kKS6BkwAj5TgjV0S+g32X9kfJNq
1frtKX8fm3TgW/mae3PtD83wMHa2JHQBdWdfDCK9UhnFEKman1b4ZxYqCU9LF/yO
+Jdi2E9c1+plW5OUNt7t4HP47RwLJ8pz1fDokMx/phN+zmAtJd6jvxEMn2AnZvsk
c6c/0EcFiHnP9MYEV3lFrRnU92yP1a7CAlf1KWbnCNkFSXZJm41hQpxeKIP8xxMb
3wRLkBNbMWIMyEK8zLdQjRBlL/c5XW+WLzMRscJ+jaMPVHhVH3o7UnkSYEs7qobd
Vja8zo5Mje+GLXzx+CFHgBL2/QHnw5rYAbIXmhexxuEhwuZKeKcUXFIT62+ieDY9
IffIih8tWyAjrfkJuUgbq2vNSTiIRYkFhNhPoGjkkXqU1a/ejHnihB90FirIaGD7
fziXLvTTxsJbpuNnKfjx8G0mtRFw+nYGRTG5wzblQUCl91iFgIgPX32avXcwUFyj
hwfux+j/QxEpB0WEW6Dq6bjOSipcmaEyNC4VTkQZZqrTXzJp7IXCqK2Q/nDjZU1t
dfoCndhBDsTXUr9Uh+WPHztFcxPDXw4+IqSw1uKY7WnWQsQGOyYRxwm763uaD+/6
z1hvAsLVwf1sRzxYBShhVy5lrGp47zGm6DaFG4euWKfs0DFdSola/QH1naZSErqg
jXCT1STDsWnu64hH5QV260FjDZZVy+YKUi3j5cV3IOgj//C/OIe8S98WbmTmaJoO
MCdFFZmc4opWRwUg4U9yhxfNwf4u6vkQUVf7zbbdF4Id8Osjj0wkNdsn6IEvYc7m
YxL2wiqJlhCv+iFGmJ6hWuGiL9iEVTNHktWMN8EstRBILxludHCYCF/vBt8+emJV
KKNVK3HhGOezkoWgqjOaW63KGI3TJJMLas2UFfmh+bUBlSpPEe9zA9zjsOrngQBe
eON1vMfZW9RIc232fNMghDsW5PXENkeIKhVrLc9EA8cqlALplC4lspG7DVXwzvjn
1f6Ssrbb/SkfMSoukAUjdJPV86wvQ9y8vKmUMyYfJCGH2nRuq4cmaeqUWZYNfvE7
r2KiUgB7ga3ZjYxJOrYHzsIkWehgr5Ybpr6ZhQcoMQFM/bNKygoz7S3aCbJVnpd/
0epAcm42mdTrrGC07QlUOds1ZPC3wv67yC/k9cz6qFocLbRNZtkh3kHTcjaFZZif
opcj7nWbUmrdyHidiAq2M2Gg91QwiNWxCzeTwEo7OdwUno5U9Nc2O5ALSvFNE74i
IMGcXMrCwyK5QBDRJLHWIetuccPOcJFcpU2hD/5UK8hyGcwy4BlBe1nLdqciAsV/
TbiPOQuUPC55NXEDEmw+KKu4O5YS0VdvW0INo1MHsON1/3b+8HktQ5S4WsBqRg2f
vwIvWGAF988UqURolgzZ8dLG16sRlF2Pq10rw+I7XXaiw32+K514+s0e2pw7aMtM
zFQYDb2PMv4cM7Qm13Ha53dw3kEH4ZcFB42w1QHSvK78AmXdC0YNRGgKRVlN5K1t
HlkfBP5B8djuUEJh0jYSCknxk4/avLkxq/k8EkGRt9WOCbledffA8yZQBlJi2HVU
r96HgbDR1o/FE0Q7mj9x+UBSyaFwbwdhFBMFCjugthSEjbh0iaSakb2rkzwmmoEb
GKNpKHqTKoAE/g3q6nKmkxyMVA3u85TT59x/4eiyCnzowexFwXE2eIS+KoRhRnIq
Ff597RKsOchYI1DTfs6ryMGPY3qFDlFkg0p3l0jh8NKhDo+XEUHYrq3BArTRS1yV
mLRARVAix8h2P1NtjRGTmiUXV51738CItrxcSfjLV0BW97w5Wym600WBwB/3WaDj
Je2XqIYm32bY7lcFhqZGfWDC58im7XW4z/HG0VpyZxJejhVA6ABt8tRPEuvkT3QM
xzX3NSn1IUO7z81a2yL/FAnkiTYg1V7gKrOw0+QzLLaM/CnCEM6cIPYQJz5vD5Gz
ER/2Q3G8ZAfownWUbpxikKH5EgtptTTW9N/U8p7pd3La6t4HNyciF46/ZzJv36xD
pPo0cL3iuVV0HsyCdJ36RkZ3Ubb+MQbT/BuRkoohb4Nwgmkoc/mOQXVwSZgBTk9N
/UG7RFQAAC4YNJ1Rfbg8BDXCV8zhD3IGYfJSmykR3rEcJGIAaoE1aqpCmrNYVtHc
L2TsBkWq1Ij1Svl9jsiF+HPHwiVSXHmnDy/FkYAzADeIDA0/zFNcCpRcN/UenEEb
vG/OM4uqZjmITaOH5kij8V+WD+iz7FuAcYLfeXbHxTX1V4IcMyLbhM4UsLN8U4JQ
EBw4yr6wqSUqXMMTj27jyeDCwJSdSolNSWFHI56QQbmygaFwwPd/xucIQypSddXN
kajs2d8ZpqOjfWKohM4HwqFhKdLbd9Z2GRdCOIUPLdkcw/K3eK89UMBbgy9vt6Hi
Qn/tyzSEigIPS8oJOISggXxUGOOkHNQts0iJf/vo38sapXk925ehLQTck5LL4VU7
pfBa3lkyMZczkz8KIYIb/iy5gC6xRF/GGXOC5oGNb8/HaAouR/4Kn7BlbN60MEb/
0F4VwJfVUQqwV7Xtb8zcXmDa8/1W3I6pOAiwAWUJDIcZ9SjNS/tASMzxn/AMbont
NydRay0BUgcgfMWh4avHW+qGJfAbXeEYHHlRC0fBBW/j2BreziHiaNpPtqXytylM
YyPd12PaAPnG4SR6XLQxexRsd7sJ6xFIDXaRsKmNk9oypVEpFUlMFygTB1flQ9N1
thMMeODOUHUgD3BzdnXIN6jVkmeJjypdTHaWtWvXeYgJbN7fWQGWwR0SDCtyJWQL
ux49RMQgm5Cad0M+HxexNAium9r3VBmFs17ZI9cGNeKj0RzMRS9UpMsmJiuLLMak
lfZVA9TRUy8ycQTBiIgqAYvLQ7Y4vrhHotePsohZJJbj4V728Wk/cFx1r5M+7Y2M
HoT/ZdvtQ4FO68aYpnKyfFn9h3j/VLBavlIjIq/mm+Ha22Zuo4kIjYFAuRiHsZXw
PJyvUvVaPb9e2yw33G+aGpu2yly5RE0NS5k+2GZ5SD/Z5NlT1CrvBokA2FGHYQMb
tAHz/1GNljuqkDA/oyMD1mUC38zf8GMTYDbQztr0PDAlTKtYRmRigKtkOxk5nMBG
Hmx5rEtUJmeNQYfpTaMLwxQmZ7OyvvS3qs0ukB5at0ipFekh4JIHyGg3sdHOehHC
xnReuFfa4gVPmOjTOdpLr+hTu2n1QwFBAEOxPvmZu9LNmAJuRoUy1JYs+WlG7sVc
+DgKB1WBORR5xnDyqIzkHZagSd9878p5Z9pGMeXiyutzCp+1JAoKwJKYY84sWhjs
ibr4q65pwCTT3alEFMzOq6WdUull0TS4upQIxUklNziwwPN8sbMLJDpEw0WSIskk
UejUyLN8cCAIKshAWEB14t3JaE0P/YlEjR9ZcDn3ks2KuFVFPt+yt8184yH0X553
K27Wv0SMNrOYIIlyJ53Wqkc0Jo1iVZN3AjxjvdyqtNYIRZW4iOeGz0BQSDbZxXiL
e1T2OfJKIrenipEynXZNMj6C0eCExP+5qCneqFpSkAUROj+FmQaksXefrxdgs3WW
Yp7Q1D/Eaus9LauarkTRx3mjaggXPR+OExCLXIwUCc0fdBRxWymW8Uv8DsOAI0E8
9AxC+qbbJnAIR+taatzT9rOlSzB0IJVWqvLKhYkHRgZ4jz+LXm2NQBkkzFbK3y0A
MiDxC1ad1j3lc7EEfEdvIpDBuZTx8WrvvuLJW/K6fhigciHGJWKJJefuyKM+km+T
tV3HKeE0WCYDzyX9nqsmLLy/Ajj9BaAIS62GLgp+vG7OKKha2M1hmfzXqE7OCopV
BMlGDQM+sDk8KeuJ+M6QsxYzmLatEcUQynvWvGtIGs0Y+/PUGVGZnFK+FCS05EwB
DUPfHr+rjXgr0VX8Cz0xVKIYEiFgH/fYVueQUkZwMrYrfd9YzGKAZdmZgar+3Db/
k5Vcyg3i2oOJVlG62Jk3OnWV1lGnr7GlCuCO+XcogHVo77urnkoz0owFVhHWtgS/
9yy7QuOqr94tbTFec6ls0mMEZNZPlk2Sz+xEWgrdo1VEvZG4jsKWnFj7ffHr8nBq
Dx1DNfxkU/Lvgc1/uQSFJYBkysEwWH/uDBixMmV5kZmeBU5nh+Jj+NsSBk2RF64S
jAQC/8ONAugVLa57qewMELy1VXOC48ySVIL+TVxz6gMOW7SwQjSHLSaVYSoFXlQU
DF/qW45aNodhrH6I/8gxyvszXYdASFbIR25rFCRcU90PHLP35ycOVQCO50i0SxEi
AZHq6wehbTkZoL2+lhb+njmO6RZbqU2UarR0qme/QeV67CxCNeAnQOZBwIKdnZo4
rwc3a6ejErrUw3/PTwUSl+JtZdbz8KGlM/dVWmLS1SyeintTlo3Xb4xUCRYPPcHH
7uf1jYXh6imddLSXUlApffMtZ1LV7nNqlLvgCiMQhKEFufmsgOS6kDvaam+Fy+ox
DgBuuyFQZJewfdwIyAU1/Ap/bd1I60Clv1sRfzSEgbtSQQgn1d7RA+JhX94JAf/v
WJEIK33aSm/Xhn7lPM14ef7PvWAv96UtF5TP8iZUVd8f9xDRHYBHxGOeqp2VowuT
Kwa5Bajh9slboOtVq6hbCqmOy0g0XkKCX7MhJA5VHZ9U+mHMp94bUm95W0P8qet7
Le2D7P0+/5njLMsiSAwnlMXC8P64AzYmlGkXvJJdL7kHlAsLReckAEt7+tJqytN9
MDl9rWlVtqx4AKciq2h7BTd1RnSHS6MfMyMPozxquvewTz+pKhBHcLttPp2B1vJB
r+C717cEGuYL9C1sCYuDtUyR+aBj3vWJVUk6CMa6eoL9p0Y/xAUmxyuTm2lFJ+dR
8/+rMaDgS9FBw56yEX+yzykm8IPFRyX5NOfFunjB3dS5elbCitdF/u6rsIj2Rgwd
Lio8P1faYmRvaeBqUPtAvK4XGLuTsaNoqX2hB5ERUlJC4H7EpCrtEkz7Ya8vKVOD
cSqugjhQioIvm+4YCNtcZOK5CRkPuP6k9ZDJA1u/Tu74/Cla76+D2s4gp6bWIgpq
3a97zIUDnajJuoO/yj2W7tsYVephwbwkFOQlgRoFVd1lRvMnAHmpJhW89ox8meYL
p7EyKSux+zLMxfQMHn4OCRxKNstLWX4BoSYLlQ454KVz8BpLZ8aNsDRa2XlXke8e
SNTTzjo7tyk/PAcOGZusKFyNlVKrSLmETd+D4E/TD0x3KP4mfnOhXdPeOC/w55DV
Ksg/djPVV/UysmGkhX1g1dkj9r1NY0lbF/sCY+lM6JbwyoWxah6s2KHcmztLdrQz
lAu10NSQTvhpkzAjU7ISrEhNkSeX7p+rusyPCyEtesE7NKIB9qFPaw8ZSqsr0p2d
uGbaWRlejJnnqjDKM2TVhABHEuoL3NeOEWxXqxX5/nCwz/Vn6yDCJsQD7R5GFjpg
tY3EPS5edT0JnAP6eQP5XW0GlXxCiO0OZEInfkw9vmjYfzqd+zi0RbJ+fIDg40E5
2dy91nbcBOJji0i0XrjDTDTUgHGdouhbm3My91JR/2ZVqx1zuZ0RydGUUzHCzO+G
CK010BLa+Fz0iYgVE8n6QVC+O1HstQ6XOpg3ITXIx4NI8JejRhk3nrXEwWj6fBw1
nAe3eVL1vR8Is5UuhPTsHKqia3MU2mvxM4qJNCuMNYZ5gsq2shZXpaAKs5Cc9nBS
TKm5bKe04T4Jlj64O7K3csptCeSftDY7kVFK6o50Kj2ZTIyrmohqRIVYgMWca+A0
8Z1yq3yZ08yWT8VXwVM619kw8OU7I7Amhd32M6+6nw8WFV7IPWsJUFZLirN4p2FQ
lIX/uVRjo+yeuxnTSyfn9NvTE9bptfrVwXtWzjLJT4QTgkyjqTGuul16z11J06gv
KAPc0H8mYTYUOcFiYUPt1wFP0igAoX0bUlPSRksIACnvlNVQFrESvTiAzbS1sUYP
J4eGZppHsVHFAvoG/fP/ZyiC1fZ+9kbe1BFErLkx01IWa6U7exb/1fIGY15jA4pv
DSQveKexP8XqIq2eiQiNreeBn1FCht/FVzvJoXyUw6K45pAOXBq9nvjTGm0fN2ep
X6oRuyppmiraYFkhlPuzlgobmtndboaI1ZcD8TQSJXdDg5chrg+w2XA+Q/Zn07h7
5AdtsakbK1EzqAJHUKYWo4bDUf9WNNCIWvhn5Zew+DNpOJdjqHX53WLubRPdAeJg
fzqd8htilt1C1955VxybPSgsunWjwa+IhLZzc0oXnklHrsVz89gQ1LM5rX7HSu73
eq2Xi3oiUZVgSTdjban70qWOu/WA7duLFt6xFy3ezOSLFALB14WxzWfGMXUudkVz
g68sXUP5iIdr5HTxXjsmQ/ghHn/ZHv6g0ECCMWy/f3kEjVcHsovYbkcBxllzDGx7
Lz/imv5T93UwzI4lIz2WmWbjz2s0eJ5aUwuhVjvNJtm89URanP/fzEMdiTqWG7Pn
fwGFF37exr/jhtTWp5XdOYJxMLqwlIg/QZhm/a0u4uXmDUsGkhejffXmEok2dpw0
9mQymjMTrIKkd6KYFFsXFkTnzWpMtwytSiXD1PoSZ/KTuWlYoANG9Mka4IiAQmdR
U6P7bW6M/cX7CSKFTcQZgQ6Hic8d3Z+gBcOTNguBWcN0rtEYUGLNk2WIjrWzS7wj
VGIdOym/a0AUF9TGc1GF35a723iwN7+d90SkOWgfsFRqarEFafHHXkgur4sjdpXP
GBQPakVyeyN1xXDj6goOeJpbUK1qQF7W3s1et1vqmHGtCCQqolICd8rYUWzBvMyl
Y9jr3pIuRLvR7HOpVT67+66PbSnx/vSfSAhP/pvG2I9Js0HHFTAZA1coUpJOGM9k
hPIYf/clRdBPsX/7LO37HdNv/IBW6rlFAJn95YYeXzZK43NcMCeSCLEfwljdH+ZF
2BmYB8C+gi7HOsq6oTd24GiF2KJ/uHmJOBDCvUt+GBbLfDdo9HWD1blgC+cbhJ8f
nlSLvtBk8BPf0MMJJjM511V6o1nX3e7TGsPM/1cAFDMMo3L66qYgR4MvU5TM0/bM
jV+sqRPq8bvMj3DPYXy1UFv92H+seoVSxGA/oInQkeE5wKE5nXruaz7VCo1PcdWR
H4QaNYsQQOHLbLW2SR2MKvw/MfGsWIDhGPmI0mkmHEBXUgen0cGmQdK29pOkAYvq
wXS/GOwy7pRcEUmaxmiJbCZyE+nkuaaJZ2i0qYS4yhGV3ZBB7v48rF/kO2m96OPl
1Gi9X+IBVvL4E8sh2QNeXyI0+UYH9ecpHRY4xbmqyNqJZxW7wAlNrellHi1YycfO
Ww4e166ufCbpc5b4uOJUPI2giMCIRlRnFYu8tUFzmtbrw4z7wgJpWSsMLY6VsoUR
C1sqF0t+mESjh2+iPP70445VbltHEQhMJ1+GizZDc5YNgjP3VHE9rV+/jJJvFfq3
IzebXsNF5p2EpIjuC7FybdloHqd1KA76EkQU2d/y02xOgZc4+NyHYVuHnnv5SKSz
CPzebhStZ01sa33uLclJzyfskgPk5vwNbKI4enFIR/+uLv+ymBY9zre9Rt+UkhW2
bFh4aHCj7dBp0zXuYyGARvzDTXthRjtfjRhT2GoRM/n9iElXnYxKmh4Gh6+DhA8z
S88k8Y+/PbdFghTvKunECsdjm2jsEIRBNz2rDPdUQyOoT9BC8mTj3mrYVprSefsb
qFy4stiXLKsZCy7DYf5NxafhtC2oE0HuuED7gKLOn2HsBwuEQa99a47wEn0lV3/r
6KsARSI+YFHTnsDs8Sk8QVVzkezVGCYsg7PxV46qbLtLC4g1LG3WjPc1Kn0VU83J
P37ebNsg3LQZQ+H5vgYmeNtdcRI6aiuey+g7qdPGfagwlRJuJZBBK+16mVbPZAGA
GBhIRURbRHiNK/7g9ayprpp0kPDE8mF7jTOD1Rj5VnXPlk4YRmgzgoPpOKnRzlYH
pjNhzInRFVIPvq+aWmCeIC49C02+Sg6jYgh05MsT7DA8NLUD93pq+HGeWkhEL09p
W0NZNJMfum/MgSTHjUQ7ItsSsMppB5FXG5tPj5cc4VLXpQ7pD08Qhqbfbnw2XVNm
X629PueBRiwjL9LCHn6DBh1YmFxe8c4KEuFRIridJwvKjz+1KfFk7OPcmZDCrz3v
bnAwdAentEcdzVW1UkqT4ZsjnuDPnylr4DTCRtzShp5zfPD8SlZH6wEWRr+Wet1V
R/McEKkvDcjZcTKM3hg6CPR4D/elm4E79QDbTAtrEkV131ukSJaDvxVu3GHWpDF+
R/7IKQP06qzQ7JPmIXv9nh1MoeDqe3Kg3QkN/p2lm7NiCV7OJphluBSfXKuYBJmi
QWeYaNvgSNGwu1L90BgpzAiPpyr/yly9pIiohYz1UF6666762KOPHd9+wxFvk6Xw
YXcJ6SKeq2Fmnb8F6odY21i9z64Oitg0Dt1EyZEAOLW3Z0SQreXphMF7TY/yHItj
XD2UCZPdNPzhMrr9lCbHlpF30Dsmg2OueS52XiHAh/Xlot0EttwukbSQAvw04rov
vY2xfVwOe4OyynDZdlWqLawUlupZiHvZGxgnCV1ashO2pqr8uRt0XY4qMmDbd1w6
Aw3dwnVmCo9BD5B7+2ypHRTegjR3wYs2spumkcooLqiv7UiHsKICXjZAG/rfLc1x
1+x4PfOAR5MnXn7qdKT8bFkGnIqT5ZmrXuB8cs8r1uP/r8FVuorzL4y/cMiK7ifI
k8K7P5YTCaobM2/RL/ELGWISI0o5EaKU14bd4EiapDAbPEfWAh3E3BMT2xu/C4LL
TGuM5sGijHU0aRvwQckmUuC2hKT9aIbS48eaN0Hzx0Wtgrgf8LoxhZ7/3whWzcG3
19ZUBEKKOHRAJQiDihF6cKd4UEl3NTGzbM+Ppc/QIlHLeX8cAuqgEGQ4w8wEcfS3
CXScL5E14HfWz5WQKVWzl8d7N65NgPhFjyJkbzGfmXgr4SS1aMgFWe66+QZhPDIZ
nLmzlD0uNSVEbO15SVG8x6IWFISz2SV3f563BgDJ4vKZ6McVyb5KB/tbwm1l0ibC
CHEebF9JC/0cI6Na/flXwMOtTXYyJDTk5pNyxB3qaxC2ui3r3ew87GmaaRQ6pfnJ
lTlJVT4vXQmi+RBFEyLKDV8pyXsn8fNGeUXftIzmimDQclpqayEe4CMTKsnhRLPA
beVCQY9oOwHEoix1Uk4YgmlYs1+svd+xmpLsnH19qF+9Vw1jQKai5UNMsEmZ1ih7
GbdThKNx/dX4U00+bJAk8X0S8DrWR0mi9BAIUpetvyCp+ew+WidyK2L4xPaz1zeQ
DJwxI8TXbn2S8/JG1Z0YdUvOErLXbsf/ooIR0FCbvje7+gLbasgStnSIFsS+9z2k
8l6gxNnPG0a3EHyCehN4RdwHMQBMeaOlehDvtuUE+92fbfu9tRzYdmiKvFLkkfcn
Fv7mnhm/BBT+6AEIh4ldoKdimGj7tN69Nr3eUgeaKcCXk4zhVShQtOsmQ2CBn0nk
qQ2f071i++3qz7yQlKfeC75e8MYw8x479Mb1QBlfRyY93xgQ2rJd/oDVWGY2pPSi
64957W3Hyg4+Gtq97I6CLRUzlDQNuwELpSdNsBdGw6HhK5D6NLxIBNRzE1ywO4kU
Vka4lWsmGUJ24ooaFahbI9W+WdGCoQmagtkl0c0LQqr2ltGFraR4f6fgaJlhYSGE
xCpS67VtSMHAaoEJZyt7ulC652G1QX2BRRt8YnHjXV3lFKkTjF4QmrhU9GXjNHvt
gBoKWZPjZfQf3P4fk5QRqeAO/YXjCwQ0BP8M5K1rsmhfvBPf3Lci+P7VtT4bKaq3
NwkcgzPdSiRHBEikbF3YoW8ZONBPZCjQlwHNCgB3FQVXW4hCpUYTW0rVxoOuU5gA
MYkPKyv7qRiPgY5dBQHnOo5B3JWE0S/RU8nSz2vra0bmATR6lHtZZmufQeIaEkjt
xzqmjBRXjuHqkorr6HoVl3V1gBvNmXCeAX+gzMsXKTWuzV9aSws7CxQ6twhQyqSE
PfbcaRealy+Gej8WkPoM2o6NSN0CS6pKiEhKL7Nl5Lw4Cuw3Zr6ayjvG8i1Uymq3
38HHA1iMGm6SDvnTJZNvtsfxqjHf3/AZjr5lF1EtibscEx2PrIFFE0d71ZGbx3Hw
chnX7CfsLscXnr8+hJMEO4YMf4cFJfxFiB4UO8NuSi94cZ9zjlSOqP90rpy0GP1W
dW+mSEi5PXM//JO5WVHQIrg0ZU+NWf6WmxQDXz+HZvG8Tm2UMM/qnQa1vJBjQBcV
j3JEsJe24O/TfiFuNKX1kWQSlkZv+RSIjWP0qof9zJlKtvTLLGd5BvDmF3GE/1qm
xo9zj3VHeWpAbBsvekQOh3w57vtngiXpw6OtL0a1+O+JouHr0SwUQp1thrM/RTLR
BZ7iFEX3LNRhjUc21XAlKmnH/Lp9pln7a/jK85BswqTUpwsrLkvotA2hL86fnqXl
FFarVHq/YoCPKS3fUgAjg6NjU9oIAK49e3GgwatZ8MbuNX14TyKFN10HELFw6dLj
bts5SbOatorxCUtdkhP6ITaffAxg+E+5fijEBoY7DHqDSE4cIVLvzsuMUUIZqc2m
Zc4AKgN2zZxmrQizr9bIx9CBLkvLpcPaAZRQol456voKZY06Rc3vh8ylbtLBnuXj
rXmYfdCohwzcW/NUQu4sR7SysX6W6uF9cNtdTmo2voa+C0YnBxbPevn1lrNdnuQg
+vwXV+64dojY4h2u9w379mJ0B7uiywGVKvQGp6tEGb2ERUw40OWTqkl6w8BIfxGL
R9NNR8UyMdKuQvg2+j4vW4z+O6jrd/eR6S+9lJjmnWTumvBfXVuia0PK9RlcnUt8
wGSixVse4IksIEyYVozJl9eojr3qavv4Uhr/Ws04FucmTNGE7EYWOBkkLPJxkRQD
XpCYUFEy27ZTR6svmFredtzB5/ocf+u+6U2gCBg0WV8vAJC7nEWILrTx6mYcT36+
p4Y6NqvDaPnrH60WuZRyJzviaeRlHIFjxu9Vf4h8MgEeFJhGC7TL7rIhOtRNbXaV
pFJxwDtiSgJao57m3H1mxbtIeStIzwRjV/j+B+QBl7wIBv0jOQGjh+MePDPKzbH6
ki3zrlJKmu8dr18GrIs4FmVqvux6BE8ERG1YSqPbZK5q5wxvwYm44/6WU2bdvSNy
Ri+4ZeJIS5KVnqgxGWKJuyfvuhE6WvsOY7ZQTdWs0aUIwihOn9hHcK4HXcFoEny7
T2BgAIPvDtIyMIoMEHx8IgP5lUZh0hGSUAPLcY2xj1rSXYhkd4xtaG7V0GQcz030
1mK8ZAeADsX9TnpvcUGkANzXM8NXbPrxTHhVxmhZDI0ZNq59s2nj6g+tvrvGLny4
ZIwa6W2smed+ZzU7e3iKdRLc6CSxzPa0TOelDgkIGRFvR/HabwMMvnqO79AOjvDK
T4faEk8JS4x8R4Q46BlcbsYpcx09ZGMCl1Qom9lAArxaGAlJJKLV/rIup8biNMHB
gJdvN7+20G3J7s1WMprUfThueOtEX9RcAgdCRPeOh7R4nxXC8vuMzYmv8ARaXvkt
qkfRRtHka+RUfmMI0tTHYU6btSs4x4915eD6yuhlmrr+MFCWifuB6PN6ugO4Qsip
Wry+VRJwqggFj3makkSQDqZvz4R1U6hIJmfajMMXU4Et3Qjs3j7Ji6+bh9dw0c/8
37AXe6Dd9mJk7Ggu6QA6RKi3q9on30T2RBx7IZ5rJGAqv+ZZ0e7hYeL/1aqR4XY0
y/JMaDXvjKdSIyImOufC2ajJ8Y4FigiW5l8vh2rqEg0mCkQ62IgFZnBHZSnfI4yc
a5OuYHsVpnznPur3zYjM9nkhFuDCAHeZnIAN432WLKEKsGq5JTxa8U6YekXOhTVc
9rget/wDM8npNbKH9OOHC17EwjJsSwYe02fjZJpzk22zLxXweX8ij+TeIz3dP+OM
ge0BUdphvfeLEJysgBZB0C83HsCG6xanN7eh3m8v81ykDjBSco49gdfBtFWIBxpK
S2+QfsQTitp32wudmsw8vqEP2BLlJqfBFFC00q9d2HjtmG9alCP8pUWofqGReB9N
C8aApdB8/7dg4ZyvdtDmr2sWiIz9j+1o+8gGZ2JmIbnTBbhM6h6gBTFdrD4DhnoB
SxNVQNqnUliHQu/eG99Fv+as/wexzosdQza2IxE8IsjtG6XkBlMVSP9dRshA0K7G
zRj2LZhKvoBLSgR2goUNJhUSzYme0pFjw8rfOqOMsQP/DV8QRPo2V4FfNnaz/BA0
H4W38N1qdTspDBXyXvIAlOFLuMq6Me23qsEL1gNbctgzT5uua1pgl9Md0JRnGETM
cbQ59S37elYHtE+oLPoUU0dpn1cQoUuhga9U3epxDzKYT3Y4/KAN2EnzfxuAHDwV
S6WFqhFTJLZM8idqjb7T7phJbqceVGOw3WrUGHqmb39JQdcejVUBYR4KCgNfbrjC
c8PQqQBjigYaMwhjcLU3FJYWy33VnFS1SWMhhNiapHs/YjnK4JHKdkPHrwCz+jng
gGw1M7FEgMW3NbQ+S2PcKps6lZVigh1YmMuu94ENUgrcofkRoKqNkktTQ06ELKPP
w2KU/aNYOCZKfDlGKbuEHscqu29urVYpMdvo5UFfiai6vZa51yTS+dp4VE1gaZVf
XCyMrMprWs7CzG34PIj99cW1VO2Bg1wj4hPgdbVGWUiYGxqCH+RglbS/lEQZAHFD
ABAwgvMPXUuz3G1oZ5wAX1UuPh7YJrR9MaH01VYOcYsCsH6xLsFieEPFAGvvaLsK
Q2+rFO+3fVQ6PlCvc9Hi5KK2HHy5hTKVmq/c6tSurfqbbDaIbVWAY3I2BKfCVWHY
rizQBB0YprnEPWq/MEe/ZVvZ3dwlgH/k2jLJp8QiHuIoeMBf7f+cpABwa5SfKE2A
tx9asftHekxfjo7vX0fv7A2I9YaVTxIgnRStOSkQTTuDeh0ES0XQsVkXSmzy4AtM
ziM2rfO8jkfVpNDGkMDtgpakaJQiz9kpWF3rSUhGzkBWHARGwI+4Zdktu18TvOoJ
9enLii3mWF9UKq93OKqs1wLBiL8eG38xdZURNqcj/vykOPl2MdUFB64I733bkRtE
0K1XKzRZSaaJZfBQmW4jH7a3QjE/LgfsjbmIR30HfvV1z5NjioV6hN+G3l8Q6r18
9fAV8N7MndKE3ilJO8EzZim1pqonOlGAPLVd8yplXPPFgHRF5x2a4s+lVzIy9wfO
ItvC6wJLDijp6xtrczd/ALCMSWXWZdIKADbQV4+r54o2E1+l5E7CB0HNI2fvm9/q
kPlo96xOb59YKu9DjvCd2apA6RvtHKIbbrjDfW33KKBRd2y1ckaVTKbA/pn46HXv
w3auxUEKVVPvGAHZS2rlxQkPiyxnhOTGNXh3DlyQN+4qhq78+lRID+VZBims8B0w
xT9b8H6qSfkBd2zklyu+vm9DnZtYL5zIy5+N/emdPOdF6sGC6AozrjdJSFOjlLAL
bDwa9WyarU7/HBcdZHPg3imctSeZPWSN1aZ3E4GJpRr/moYvoyKehIJstvvgI3Tg
cuKB85MoYeHJZ6Xu6EaM9dtF8jUBtBvUhtxYFtxIZpGGk2XtBCJeMw8dXByUowQl
7UBseQCX9O4WKEFV7aXk4ps02dT7eRyv5NZwrHlkeXqwlSTkgS0KnKIFMtJGG39w
v1LdE0jl2TCEbXMVZnp2GlAHjGS8YKVp1nepkI0OFtiDTmA/CBxWkCEd8Plzt1Ja
frff3OzqJvkywySvLk19/uv9xsRSaRuOProjZ91pmmpygfRIyH/pS5oCIr8nOjGS
rzlMfuTRaqOGhUvkuEbW18IwwlN4mE2f/3GuPaJ0r/sXpq597lk878yi11+B6Ccv
imSHDvARtINUMdxxvqyqG7+sJzRutjqIJKjPVa99dwmygJG7NmAKLFyp0klFjZoa
Qzs1g4lnux71m8AGw44semKeX40EC1hcj7SQh/XkwzzZdI5xFgiuL3axTsDKEYTa
pZxmNyvdAEMtph8udKhUapb+eaFGSWPwUTELBlDcSNozx8TzHz11YcrecMizlgiV
axHxt1DEwM7K6+Nbi0Bn3vVy1HqCK+CYtx1I7gaBHTnNtZrwqJHcgzCIFJqahbfd
icWjvn22TaKG8vndjwVWxdLmkntGV5SZ5+OiZ8gyDnf7tgWxV4tguIqlwAdF8ZvP
otm87HrFLAMqPYEuG2zU2LOJyav9lc2rusC969YtYSn0EgQX+aPoTwAFy1QOHklE
pD6L8bAjXwNl5SBjyZZVBGvZOHuNe90HemsKsuDS8B0DhQANfVsYeFhY2HCzClpr
5De2dP/2JRKvjMXBmokcR89jMDxKT1PWnXA2RQ/7zY0QQ0h1jDG01EoK5cSW/ySL
Matt3TPhyhLWWN/2XQnYMMy358R2Dngh2azB8AO4d68VYn5GET0YXTYgl5AsrKfl
pHjdy6A3yQnV05COv1tXSG06NB7np8OA+tb9m4ZHFUFV2LTAiaGHRP4UBARKoF/L
6y1Y16oD2d4kLxQh8dU4MyIapbDX5BSAEIvwraZ465rjeWy3rQ6TaPpj78HFjGcC
wUgC+jhBl6tjf44CN3Bd/OSlipM1UDmMCI4xaqLY0MVzxlD7LFW5HADD4AoIWTFF
PvlAXrSXtU6rADVnLVW8033qYRAWMHCktrajopBkDXZccvq+VJ/kPNduaQ7TL/kD
x6C+MK3aP4ionuojoox6c6zZysDRgmfqeoQI2ptbFjXEnhrTlhT71v+HV6RWX+mY
l+hErvWAouEesYX2HvY0A41p/AK3PIO2kVkGZUekRMR4S0Zj5+JiOPotIFUFcNjO
w6Lv0dpYABPShI683VTb+4DHZN5SiypItnKggs6d18jIvt2eMg64b/oaEM/Ssfq9
6WEQgh77JKCmJDSLwMBH9j78JM77esI9A0CMERXZSHhSrwb+uslrLGGaygj+nEl3
7PklyouUOoR8yoDeZpljC1H0J65J7Kk5VP7ZtENhpafPrrQscCB4W5NEWFL9+7eY
H7eJNGdyHBdh1ylYPmL8RVi7bHbOdq2t+xsmg4L7qqK9VfsaxmI9KXIYLMV68elq
gzJaVkEfsa2weUmiYn5giV7eCexZVrzPnAR3Ij5rnMDR25LFv/KWTWQ1BNJrsA7r
IOeDlZa6xHx2Pxf4nTiEg4MVLRUpa0R+t7NVgUTTddLCZnHHOWuJ4s9paRMsPBs8
g6zymitfxairBYoUaRJrVM0tPSBJryzML26xShvmRoJMzFgMvjJT820un7qUjzlq
hmhTTE2orjsLBeJN0xjDYP26sCaBmmj4gMY2JwnSFs48OAEeA3htqZnDr4W3KJR2
CYlPkR0xtbPI6w7Q7oNI7/Dfv4amjPjfDxruVTO+4yCgdu7s9iVs3fa2rmia0gbl
zm0AlERCCW+DGWDpn+cqh/WUIaVuHMhovQivv1OHBEbK8CLYr9OUzAQU5E5a9bR5
1BKDiVjS1RmQs5xJ7KVwwagAYIPmGdan+6F2h7pMEAxClIm7OWrO09q5aRFO9YUA
BaKTEKaO2KKLxz4aSiNS/inwX6+me4XvCQp3Sl7X5+35zggK7XBr5bOKmZ6Nbwcs
cNMOe126ywPcphoJ+JZ4usme4nc7Qn1U4YPIep1zRgduawfuGVBhSJIr4J6KcgIg
EYl/fvPzzbB/pcR3KBs9zmIaK4K1HfWZ87sfONrUWFc8QH5yb1xija2MvYwyhvTJ
2078Dst8GeM5taswvjUSucD+EOZZ4iyVb1XoRsLrcqcaZkBH6xU+GPHA4ApBHF6A
f3UJDlibwT+zGxyfUIbKgRHp8tjMRKG7VAwh+kv0zN1g6dJHb+R44YmLXbgnK1Av
66X4fggFJbPN/QzUQwNrEUDPZRqXkHy5NdllkhRqRlW1Ys0tL08Hd23VgPRZ/tEC
aE/pZVnSmoUAUXSIBZUJvsrFXPUw8DhjXMB3FO3ncAte1QK8xa6YGGsvUZO/4HXc
kkSdlJUqDoB9TN6N/omGMHhYdnX6C6NigenhtXfo+IQPW57iUrZXhtTjvOhQve/g
DQWViOxedV9dNrzd/c8Dcfu+zqM6GliMxxoFsLNRbL9a2vQJaHKnGcWzB/l42NEu
6RUAtrZGRwFlSApBCDK2LdRqNGJzaUvOC/n5qji2PYjaCDga6EGMYjZY2oSWQGxC
JzxTW6P2h/XenAxVReAsL0JN/RL0l3xfcq0y7gliTpB4SpVYXJ1rM25/NZXiTvsX
TgdRybxPEwzrF66PKYU355maDD/YBMsQtpEwJUljRpsYJNCOjaLpwoCKHJXZXsDJ
jWbbNNZ2A+gi+nU+yj0+O9eBvf9g1mvGni/rtLECYEgUcudROjlQwVjEjuFmkePO
7oqXs3WQPQ0duMSaQPxje4qTWb3cEXIONRRghs1lNjhLZY4nKrcN/DIhAYVpNu4t
sN4lZW6FOMs4r6FHIVdmCXWolFW5Kg/n6wXg4mRgxAzmCMWgXX6YRB85rqdVnKsG
+gFb7KuuI5K5CW/efcHIWt2filhbtxCxTCPA8+RUN//wuBdQf+qSSC2qMgN6k+Ao
pjc6KBzJ09JhSR1A/fBD6aV2HN9YeBJVQsEiJqD0OIUcVI0l+OZFpUOJoU3yPpoq
24Smce5dkbKBv4GyZpiFVCN2/EUqlXqjmA2Wcku7Rf8xWxkkXOccV8HzltlCA6CJ
WQpVAwM/SrvdXUx7nxObXH9PveVnDtB/Mx3F10VYhk3N/wmW84tAfqrcTHcyT9/k
895YS9s5h9BDti1dI4hdc+qKjlMKU0BHmAC223Ih29I8xSzGgrhD/4aiXVAzpJX9
OOKPmavcQTyl9Rp4oq4xlwRy9OyFC5JmWkA8NMYKa8HcG6LzIQEFqXZ8pN4jo8pZ
6PNl7Ez0n6vaxFY8/jVVQBBC1IGskGt/APPZjPzjwX18RmbRplHFIdwQ9oOYCono
MDKVYYZPwLCma6iyQhNRI3QMlxfJ62csuF9c/42s3X7bN9xU7rL5B2/LC6D0z175
nNbGgiLMU42t0NRRMk+sZyOEDNFI6A4RknNpGQdMjjocSmCtgZrv1XOzpq7JeUWT
lOybeBBKhLg3nXLLaDh7m7htUJEJO53Al703jPVxKY2J+n/EOGnapQdp52VUiogc
8/w4c1FphEEs15wnnnhvayJFAdHn68eoyqrFPKgpqDPr3I/75ChKIlj+DghWRLUd
cvbhbGJIgjVqdOUNYJGlG3ws8+2R7dIsBOzvuT43Tt7U07RiEIsGjQoD1Bwtajsd
PPGXgOf7Gq8OlEPaWjUBG+LvdjDHJgqMead2Pf4b6p44t0cSjOIJFDVh40tK4Mrw
7lO6tN095kFnUE5fC4DA9E3XL0LVXknlDgp85jsQGlI1K6QytjWnnhwf0nPEQwb0
OKq6cmA6XeWYlrSumgE0A89laEipSFNl5pUroJdHT+M6u4Die0NaSIKQ7vjnYg9P
SWPgy4gvh7Wpn9PNgXvICif2gKqi+fpiiSgHr9OxZp4XPk8KJmFuljQpssk42dAW
lypiFHAZEn2MwMKiIMnfqr2kQqC48py4P5X8+HB66H7saY8wdFS0R3rztv37p/Cs
0fHJPO0Qj5CFePv2fKyZv75cOr8a4Hg8Lz4Ql6gp476JBaPhf9paxofl+6G3QQX4
+yu+2Nsr7Ux3ukaMg/9A+Zhg2ddNnMdUe7+KvhZ8eJGOWL8ENpW8emCho50x8jXo
/ZV0E1+DObK2gp98D8CTt4ZB5H9+QGWs2JOB+TF6SQj6vLOxHcNjuio8biHqYQmy
p6kVhwjs02yzJ5+LaSGJZr9caYsFt+g0iGCkYX/k4DwxukMgtRJdShK8jHqok0NA
Guk8+BlDyrxu0Fh8S+0MJBBe9hrrL17mHs1JaYb960kuUx4sVR6nuiab7avo8cLT
73Psh67/qOGdC3iMy+qYH1bpz5G9ZkW9Gao4Q0iY6SS8vN6ulJcqgRoBlj62lWPL
ccCT5ZbJuFxYAz1KMdjgB8Z1rIDI3qCbuJoAht0LSq6UH8LS3V7jW3tFftBQgg3d
pFRUc5dj4aV+/ArVDvSEPo4ko42QPoVZej7Wnoek1WDr1CZzLnEEkj5icqoJox+R
y2JQqOa92rTOdewRyeQISTiXMpFTq6JxgVPSQYdqL6VZh8YLsq2HJDSjkay5Wjr4
L6GO02Hj9443EAhhwBESEmBimg7R1CJwwuowMhDEJdsrPaBUABuoEPeU78v5IVWL
m3vj9WcRP4ZL2pVHISBsNKyQISZVPVAPGQlvY+p+SoLlIBJ13nAxoZxC9Eb4nkYt
uOPtxwARf3AaOgLkAjx+NsNqGJR+pf7WBsjFr/m4e5k7vFFM9b1KvFanDUkY40j7
Qmjbpl3dDlzTQkhP3dPPMFcuhU2E2nCNw+bXIelHoX4atW5QiA9GyXxBxS+tRnp+
MjOWUzzIUK9Cf071W5QtEKoYTNoumC/30yZZsGJPy5K8UbTyW72QgeYZHU4cTZbO
/VaX1QWyEmNo99+y16VIUeMEIznAvxTewTcQdzB7ZW2FjfJIAYA+PgsYxrfSUFYe
phf4PpYv9rRs8y57+BSomUnNBiuGA9csN/fIET20Zs7wbnLxxt+joKmVkPLu04p5
MDMeVxnLjAoKndIS49uAR4EuyxL6VcV/FXtLsJO6RUiCn9DCyG56vks6Jaq+QOLD
dGJwR7btHPuHWRvYCWdvhD3qWXr8AtEsj9brXvT4Ct4j4/crsiLeGVFHREU/p3M/
iSHiiQbG4h2QrdYowQqn7srgz81eV+ac6Teeu/s9xmDnpHVkkaN0dHFTlUyEO+tL
sLy6Xn6pljU0k4xREi6UUnIPVus3iPEvZDb7yRzCl96FARUdPFOFJrcXktuSZ1RA
X5tKwuRt9uk8ykSaD3O6t1H45lwTrQp2NlGt5bkIYkh+/JEip8p/jB6wgy3YuZb8
4ObSovWlQNE2cE25tOVhG4YXDpS1gp1ohOWzxtu7Q4a8pTpS1rhf4lZUPd0Uflsw
9ybMXXjrQ8BTcZjSp2YvFcXCbSdLmYx9qC3p/agp/pogpMOYDsK7NjQWWH8Y0sC5
9IrbH3PX0Lsv3WPxYlJd8ho6KZcfUnHPwdT4797lRSre+Ibd8UiW4j1Z5C5jYq9c
U3j4KaRsV8w7Jds/gaQ3uLNGnOIibfLRDPq7FfCNg/3HLOz9cLc5Spr9WgCI8d1n
wRCmsmtTW3QgGYQkCneuSRypPpM4SaefcYyUqiGaKg/lB8Wz6cGLblU7/TEmHkc5
eO3NkqCbM6eae+feL7jWMXD8taZU42Zf95EFmKY57EBflXyf4Fk0zeX98WBGTKL2
27BsHcBzX3sZnODH6eDj/SuLz96NllraRiTE8dn2//VijDuCZGywTXQ7qwbiRbUF
1n7Dc1HxA/rNZrdbc45HGd8hQpBm4YP8VJ+D4gpFc9s/W7G2TV50YVsoUtvx/oD1
spJtvaxeEXPTBUOdHfOmkqCeeedaP0NL4rzfrGZ/8zpG4szyE52GqXFMyeNEHfkD
GATjGzb5DSv+BIlqY/RA4C+yqiExSt2//4Y9+0nREQMbVlKEwH9fB50Y9D5pKVI+
3zppVNtuKQd25Exe1uX9QteUek0WR1MtUIU0DDH64vCTd94JNzQZ6fAbm94Wdwm/
x68rjSh+TTq5By1/71aYUWdnSVpETWsnw++WKVUNJtaliiBmr1B2bQTxheMbC8de
qX/h/z0XkwhJ1P55Ke82p7IiKLB2k+XGuX5rf7gxNhu+2GnqBsEpb3uQGOh+/tVV
qa9xO5JRIlrr/Pey/FddM0PINHa8EPkDIiBVPhydOcOzqVV8AmToBUQLDfYImRG8
lKLesgfhzDuP7p8Ki2j/6DfRXIkrJsECMbQoTN7YWeUTnw4/XpTJ5/xXFeCRRHld
vaW4DPGtwXt2J5POIu/Q0mAJNiX6CjwwOxAOQxMMcmYhlM/+vUXeWdGvdlL7axS8
tUwb5+9lycKRqixcpDKgyG5ebIbOk9KQOK0bdbnNgf/CD8zAlclBQtFoaT0n4pA+
JHum899rB1VAwKTlShPs/E/wFmzOoKTr4cP65lv2R8c+ixIIut7udThV4vV6RPHg
Usb824eoqI0bT2q6spnVRqajbCNfW0mtEXFwBgI0g76VWgK08gh1dhr7kH7kCNCB
xvIkkV36/8B0uDGEkoYOjf2+FJD4GDmVGgmVDGBPv6kmg/qlc+bPBnfcUjqk/SFb
TXheOXBMYME7gvsFR4OCQvp9pz/ZfEUIPcjmRG9pKvsacBaBvuubdqeuJl3uC6o8
MqbNeuojDq50WS0NIPbZMFSMJtVnbmItkax5bBQMJdp3BzsovADgg7vR39ZHk1v4
fhOIju2zAnRZl/bNwj1mzL7Btc3eSTEJeGq2jWNQipdi+ZGbPeMUVF2UHLuePqRw
2euCBxwpCFXTV5s7Z6Ndb+42pudFQcnQIjTAqefPgl+fKWPVoaH7dwQ3psY8M6SI
HGmxDT4xcRUGdnyDIC42iqB5+Xz8P3x3fcPbIkCDF6gBr4YiBSSR0MB8MkldIJUL
TTdxMhYUD2wKdESFYrM25Bla754zKREO5wwLSww3pQXKqWavdMOiRVPefqP99noa
N5g64lHS6LF46DygnEekzwLwTENoSdYqx0tY/5UEXBZUzOQD3IafkSHMruJhn7Pu
mWGgVZvGpaV6zBjclvua+kB67i91PJ+MolgrJ3kxItcu8NbPyi+I6Y2qrdwSCm7Z
EPKSCF+bnU0gvWlqU6a+oxeMTf50eC2vYeW0ctr44zIuQuk8PDFU8hlTA1nWYqPH
iXiruk+1q7qwfUvKadSbGyUo1Kp5aZA+TzN6UVuifsVrTiHg/8Jh5lexYuykgqUO
3EJfuTNLpQ5cVUV6WVq2x1XIZztiY5beAq0ayGfEdjSNVUGNjuV1vZYXOWvabvVk
UE7UtJhEMnvoAivhzdBoC7XWfcqGuwRSD8uh4+DST1bdDMflCQdvLAltkt4KonXL
tfajxb/Gh9hl8TpFCibAh3LToNhXmsZCRlGUnUjtcFn/MoapqLXIPhya0m3i0PXA
4m1COZPNChccXlMV1+wJ/XcUg/AFz3xOG5XzPrzJbTA+YxGCt1hnEKdRYLtUdgI1
iPcwOFIGiiztjgPwLOPR0wVM78akaSfjvoO5kYnou0RPvwxDvIO9nyeKDJ+cKdsB
JjY9qxAx53zpl6TFD1aYFT9UgCGynQYfo6uJCSn2AGjVX6A16uyV415LE4pd+URF
9f9l/pAHkt601vRq3CT/iL0sFPkqasSAoXDCyXmyTXw/ByZXPmg1bDdgdrBvFpi6
jE+znHEaI1EIBOjG15JCwZQIFtzYYitiGC4OBH5vb0xb9oe/Lx/dtlS0Y5uJqCpx
Am7haxftL5o0oivRC6tfnKkjY70d/z5XxqQsImHzvIrxIsWMgynlD5sTh6KyzTMH
UpWagX+aSWFA1bid3rRZyH3k/PXWFW3L7OdMemgXign/lChLVVBXHmsO4Siz2qTN
8Mw+M4gyZVZ0W/ztFQymisHQHd8lxtCa+5etKQ68qYegIKfYyd4K2pgMnxAbJ/DN
gDusEOAeiuWgSmeE4VXytI9q7xp2ck4whZYnak6lw3IbkUCyPby8JYucxINoe1wE
jGy2r7pHcF/rWj6iNyapytRwJAdojj2aKgtIzkDxrAuXW0VN+2hBZtDYmpD8j3Ti
PwWzv2/s9tTeYYFCtcD7RAJTlVD8w3GZoUgctDiWK3XP1lIjNXPGztpbK8tyK6pa
zMBJW3w8vZ7sGzutwuf8VbcJVsrd0N7k+9lW0xrvnhESFCMM9RoQaWTTYCXLLaBF
xIM8wNEdCXjqE4JRVF3uHhF3DSNx0fXmkIC4+EiXW6azCbOHM6nlGSU6QY+B1q0N
+P/dmX9co5QKriJR8WnKfbjWyjN4forafVNemkkcFBJAuAHP+uaxZ6HSuQVCGEAr
2IRdFw0bcoX60RJAnxsp8zIy7MockNnKpUoC4u73FWYOKB41yoQalLGIuZoPQnLc
wkVX2RsdlWhSEQEW3bysUUkU7jetcPeMNi7VJKJxqQmbB2IKZixGZ6396o6cByWs
K2ZLuijIzEWffgVwrg86HTQc/W05ccuL3mLDyjU6W+a/5skM/sijkJ6dKvd2Qjzi
g7ai6VK1TMZMP/u98fVtL0lT2v67x4lKJDO3FQVE8zcbHTRJoSf1KmNtSYgWrIn1
NgWsX+FQb+TJ3QsE/B6h8lq7Wqf3HM679ebFXim1TQbH5m5wUv5tgo+1g98Bm4Oh
fOf4JWTyUZ9aJR4SKHv868DDBwQ85TWjKuGKE1p1n9vg18Czk60ik2yY/8BAOhjh
9YQ1MpJme8imA2Hl+gkw5m/JlF1QNhtq9/vi+Jpn00MIMd5VUJRfZpiapEYP3nrz
5XAuZ3MNjoX5Wif8c8N7r7bddO8/8BreXOC2ly4KvDWVq0KiJdj0Md0cPbFLdJGo
cXPiq3rlzpDQsQTKX176ykXkLC1F74UKwJ+Pozzy11N3h8ZoIF1t6z4qZMS6o7tc
xraRO3JoVr54+5+dCR8EDg+MqZohlEdlEVL4slLyG6Xc7KyAkgt4R+InWhaQc+BE
ENQeBaiIlLUhGcsdXp9zy9mZ86pvCoqDLWmnLKt4dxdB6a6cWDLR+NySEjN2Ylvz
bKPriJHUaNqLTSewxbOczBbzAvVWElIo1ZS3fufMRzg7yO8+5zjA4JPraU6VRsw2
8qntf9DicLMo8R2rjiVuU0fpGkET8Q65RGVHYRDsnKhPWyWqsFUS3aByh7b9Y4Q5
WylKkHV/83V4VH/ligNoUhoToMzC+UDS3CAJZTgbu/87hHRc4ZRnXA/L3ojpQBU0
eMdI5C8fveVcyn59EqMSVhe0gM+p5SNjBVNofyXtJRcff7gNIzbljwHByDYk4CY2
Yr8HJSTZOtOQFxLPz9uKpGs9FLwGBFsOFj9s+wmEmSQfreqDfGlpPCYaL6dTRS+V
cWn/+3UJLVCjTiSViE0grKDmaFObbQrjslfchyjPAOp0XJ3+DaALD5YhmAta1lRy
BidxsZ1RKvroq/+dBltDolNE9Nhyxqd9ZsZsQE//FOgIFSbk6v5D/jJqNZ6WVrON
c76vnL70A1euUMikubPUOvF/z23VxiMdomu1a0XiM7eWARZSgwLVUVxJfbcUCMcr
/6thIH556K6VQm4AdIhgJVwTQ8wgXWF4gwqdU/BvgbqDLfiIoZpDc88+F+AvqBkO
b+Jtbga0mUZNgDPVYlVB80EumuRTRaAQRavyXVWwFnYnOX8zr41lfrTygO044aFn
9I4W3sFrwyLVolTv+GQOr+1PL/+Ccoepg9SR4TlTSmly3VYTd5SGmg6mmurbF3fK
V89CofgLQDYEH/jFtC+ujIVdbzWv50Yh5RxSxoDHjpodFEuhV47mYdc0Zr2kGwk4
P5VSY92pqmCIyIJO2Qre6X7+bJDdNZ2H+X37YNdw5BXPqeTg4x1aQYEzDlbHLUuX
IgXEzgrmTsMQvzKn1ifxf+fsAXb6ef70hadZuFIbfsSykxariQWIeaP4oIMHDWJh
DP9RAwIFDu4lK/pxdMVfVZG22VWMJOdqaFzb6z2SyZZDiQxkTKOQ6BeB7KOgqjX8
XkF0yhW/nnTPjbQq56Y6TnVq7MlbBtFV+hrpeKFTnDZNh0O6Wrtx8pX9Oh1eckLI
Yux6CwqL478EuL6AkWUW2/oCd9rcRYxuwch5/cYQQ/IzyocD8xzQqpgC63FqoGy4
CMoiGrH4YudqD1aeM/ZGxfEHS68sMRBeCo1D9nDkh9QLppcojMjZ1Vncc8k0OV8/
6YCYnYwHWI/MUQ000DIjJQhu7ydqSkij9sTBaZHmO+ym6BlkI5bzxA24RxUNIiD+
BYAI0QW4Z+IMfp2rSrzWumZB0VvQWCuA7J4tTD4WhU5y2YjVleM69yP3G4Gr3r9Z
XuPaGFIQGz7TM1eT0NaAhkmrzCfI99e3JDeOS0z2xVvr/wIZdmw2ohh38JjP0VwU
YfYvrYE4hYEbcdWEjTreIT5lGCJoB2VuLPwBsPA+lkuWjDw8YYjh6c0OsM/QlcFn
HbkC+9haSLQnAoQrV70Q1NeB4jUCs7Xr4WWmF1FS3Zp3KrFISfs/Qw2KkYdB9DE8
/BAs3j0VSHHsHjSd8Ex+7BnvMoryCEUcodBCZCb64bAwLa4l7jxB77Tt+v1xR2Yd
ogR9K2kfR9pTvBv0H3DmngVUxh7FnDPPJd5d4mDjtyEZakYHgFn1kv6shbsVikGg
p75JlH7y95TjXH3A5lHw3NIsTkSEs5GOK7rWXavXs92Yf3RigeiBfSM4tUZzgDz7
7Fc2By0ajXx9TGpaUbUVcqCFhGhMzT3Xrq7RDNxkdeO0oCO2ns4TSxmxlF5qn/uc
EIxLCxzbY/Yt0lW2nGxwruXVICzj8/jfxXa84bCg8EnSLOMPj9YKEwJzVhlECqsP
Q23MWJPR1uji9BkK5Cw4uNFun5RhDRfvZpu78QdDsupWEUkImNEofiiYQuIOCfz4
5jIpPzqyFwQ/LMNgQ5XoGRiAN5Nx4xExcJqW/Q7atGFP/Ye4kr+4V1amKdTEsymO
oGMEHWNnJnuc8tssCzlCyLC/EfOM3Dx8fDsc0dISrLQKaCYIitrdRGCjMFBxpQeX
IRRSFKjQa1vddK7fJRxl2P0tRFLv66LxJ3FIJeo9h0wVouY4JvMv9IAXF8qQXgv2
GuzJOfTpFfB/DHa8Y3iHKYaQhuW1syc3Qc2ThqWgdWwTsCqON+79ENmjkuFkRgMM
azRXQ8D4f/qFk01Xsd1WGARAaP9MZnyavmsopwgGJlQDy3QLz+lJZyz21MlOBoII
S/2Py2SAvZ4/JODrZLaX8YexpSAR60n97AZc6JSnml/ULw2cCQPFSQJ0Eb8uSCRJ
+MKNRujccg4fR86RImvbxoxQyH4g7wBEfnXoCjvLfNqHBJYqm9R+ILwSmu8cP/yt
vQVSsodQLKE1dtbQJMWgMAOUBAwAx1ort9RkAFMeUQsItSVDcDUEOjLQJvjZz0IU
XrTvaG4xzZq7Rje89Lvl++p0H3kBBFCpesjR+7H7ugi3SW1q/42YAe6X25ohJB5I
FcY4QEq4SBla8qJxXYLAXXfhkdwtwzv5Io529eGOYwbrg0NwhcszQgr/tQMtQsQI
3l2vJXRG3skGQo3De9q7AaLHVBX7ZrJJbgZeiLW3C65X2Jb20ZYkf2O9Eg2jxFHn
/Y4lR6dYcK4EaSBXuvvTPY9bvbYrqsB2VTOJB2gnz0tplXIFXh4M3AffRrNTRaD6
pRoK1BCYPNoufS2VcHBe6Jk7DRVkvsHI2J8ofK3Zdy03a1i3/bwb/vsOwKnqhVaY
0o6GHF3y0hCZAPHAwUWDhAWpLBjtKj6RxF86cfWyMv/F6xq9PThGz2rwLb5Q+aOp
9rdKuLv5QiDcbyB8N12KDLmXfkuZAa3WxGAvK4j4hGFZiTvNmCL/aMT8ZlqDzrbh
UXzRUUHZJyZRTRNShxhswZyL46coktKzSkFzmMShLJjteOSfCD6hD7ELlHDqVo2e
sOthOPsFTH8SRaV6KkGHcGIeG+iuaGXIoKO2/smWJ/xPcR6uyRjqYu5jpk/A6Xvc
x18vJ2hyO7+ndtDRmPM/0h6VtvLG14UWs4r1cGIrkRRdFwCGAgZ7GWOXuoDxSUAf
D78MFMbO62oWbH40aT3ELkdGTqFel1UE7IrRSHNFJhF0hWiOCF4MbYFx8iteGJLx
MOwtkQr0bYQmuOut8EDsl8mt9UmZJYUXeAFcoSxqMM2Z/CEtcpZnhgadrD8TXY4s
BjL7i63OJSoy2NoSK/c7kpAqMijPDDu6udC4T08VeA87DduoPA0IT8PCkL2+l4oe
QaPNbIXf84GJeSsEZNk8m0X1ar5dGFKFKHy/Q7ehE39v7bzcBrmibiyIoOybxGic
M/NO9QSeyww4dtZDPknjeuncs2qPxBvbdQgJipcPyfq/nnuoBTf9x1uJPxmLb/fU
8fJNCKeR5/iy6fXLXgcnFbQxE6SMnN0o67PGlPyU3tvyjVp6m95pFJXvsgdV4UZq
pPn+rpRoExLFpOe4sH5G450TmSnzfiGTConOnc428TZnMIWZ6W2IcLBof32X4zwM
kbGJ8d+qUnDGBRp+qbGsIYiUD9Zls63D55EZP0NCkaaECi0CqIKxIUgn9zHDjkL0
VZChZRVPNv8JlZgUwfMReoJrvvvLlmKghSKuFwt2FkgEDei1AIgYMRznL9Xz4wVO
bbVqVNK40fe3CCz2y2m9YqGj53MNWGSV4qsYgNbY/4uvMwKEEahBb6uiLh8Hmla5
OGT7+kG4gVO2fUa4+aXDRcdY6yp0ck1NckDhvF5Xg9h7y6+Jl7zIgHZ5pBSWuFAd
4skkUKIFSYNXpQZC6fXHUpwPLNXNmP6osuZYxQeXyZXOXIIJt9d+OiKAzjBK7J74
/BHB7pqys1zVAGHip4rMykonO6KexfgnUcwLSwU8GxoopefXKZS9ZnPqMagHqPC3
aTFe6zzyBwr3HqM1JBDq77XIqjIjs66o0hwfgWvOE0l63y3yN95LZ8RvIOlL/hGH
ccPIBMhm5EBbj0ol4oWMJq7aynizuIzH7+bnrMyRsssapfr2ao5b8lTe37bR/Mwy
zC+0OVJMa2qgyX4OaFJmpx4KHHPYx4YM2qQxMynfEIWlCO0sDujimN7PVPTMZKVa
chUGH0Jpgkof6s+/mSi+j/h7gz6icc72TqgV/x84pONnzWwBJCktirhTqUzkAjbo
gvClBEQHWxvOqBWQdDmtxgtECToIEBhjs/+Y5KtQw6Gbc1F3e1Z+lOAsyKc1HPZ1
4tQ8PQo/B+C+4WYD2lJY9Ecs4X0wEt0QzCENYJWl+rP9TlHYN2WJqAlnSxKhtgqd
w6vGL8I/gZqMeGranuAoioqwiyoxt0JUXgUSL97cxja00TDKKxnYwlpj18JOJL4t
iQUan0Z4rE6FT+VtImlpS9K4Hg7VjsfArinKhkrc+18coXqIQlNyJDzqi+6wAzPC
VbkgXchmYljcu3IDzQknWLjf31jkyH0tpAfOvisT7/3Hs4o5zADRcNVI8s0tNY6e
MHy1Xi96UH5Bj5jRSPqQmOu2ZGsVNx3kJPyy9VIx+vkG34U3Tgn+NIoBrOScJ3Zz
zQCoC5rXX5ghjDkAdk9IIikgdyT4Pej3US6GW5aP2cr62YL4x0Y15ZWctlTN6A0u
sHetK7+gQFExLrv3SRM21Eyf2RQOf94Li3lmptAg2H/rBi/s5qr1KP2VQ8EeMDrM
gCZBmOb8gdbH8lYZB8OAguhzojUyYn8P/iGIppceXwJxb7bWQpk1cOeUp8GFU/AY
22Tm5ZCNk9RsQFa39XVKEzssgVeK2RV9Y/RTDuzBU16R/yA1YqcH0FYnO31wvIAJ
g1T+KPa+DVTS8Uj/rhzBKtHyXC0F2qkJqhCMqUm+zkR/y+kua7Isrg0frcuvs/yh
/nAfRPB7lGnAQk1O83WhU7MOl00brmze+vMUftkytLTMiISbspMEY4KCzRDmA7gY
7x/MLR5zdFJa6xfHJjMuCWXt01pjldRDqCC1dtixeCRlikdCjaAgafRQUO+OZR7l
4iQ9HW35skmJsM3cK+DucIDmGE8qR0T/Vkii/jzmVJQtiGw0/hTkhCyZEzBBAbgW
hoMUICJiy3+zFdJTY7V4OMbN/XbenAQ3ZJIPJ5bl0zh8EY72oRFoPTQSOJis4ii3
n/WLSHWIaRbywJkpmoQHXNQiR3Mc9d3X3f+IqMtNYuUIrLcZR6UM9iUWiyUcwul4
Puo43o7xvpEiQjQXEl33dZkuPQ8nTOYbDnm5+XHmO6EQX4Y+UMFrMXNx18dH5+GV
2uv46eJNlHK9g6MdD0v4/M7+Z1P5r8sPsdKe6LD1W0Uq/uzzDRUEOt9MkfBTJOjA
+EaqtE5IGkYcWzYAUWYXoiUaWZvQf0AzDcdq+Sq/v0h9ut9WjvgEpj2QcBBGam7k
BlEh2srvTygtO/4oJLZ+o28VzBdtlTuNx+N5R7wF+iHx7JjXr1KzugFV8hhwzpcd
4Vw2Rwns5PGoPiksb1Xo/RLErc1TqAJY431Vf+KEzqI1GffCwhAv44C9Avt5Qdip
prYcDQsfjrkQR45bYSvpKhbzc+pQ8h+inlKfHvwx3PuGUaN8GiYBFSNmJ5ngPEV4
RSz0zKuAMk/Ri8mxsnkFq7M6QpBV84xvu32jMTJ1i+0gM6O5RZTYiXXqr18yomtS
QYClJq7T0yzJ3Agxd6d1O+KCa30em7JSA2h4JKs+K6f1I9wfL2XwONNoduMcBQqn
uP0yI3creHIWFrpcUm3F87NlW3mYfHIV0TWftJCv2xdn/znPz/ZGmkVILW3p+OQ2
u0/d8wJKumXObxPqnF6R8O8iSqhc3Vao6DqHlKdcY/surSzmZb815kMofLUMzSgV
wuiqYy0RdoTTWq9P/axpFli1jqkucPWe7/w5RGN1le4oT1f+Ui8IUj+tWcTWlMl5
WPr7CK67U2FI5BQEjuj27VNGzpeSxoukpAvb/5OurzQnhGCm7WUJM+7ykrkNVSS2
9oUrct4pEYwzwAaaONIDoFRTvuSfvDgiOFcTlYlvsGEIIdenfyS7VD3Fo7YSgb4n
w+3PegFMF+4So7VJrc5TBPcKMlf8IFENZjUYCmam4DuYT2APwW0F5r2SBF77p0nT
fEikL6WG5TYkRoS3H2VL2oqXOJRrW0zUt7SdNZjFfTRLVBHs+bG8VyDYPqPYKVL7
9/wYAVzEgj3RmlBBRUR+oQoGFjTM+t0eNKQ2nrBTXImMNdyw0WHJ+qYkKRKHj+AM
dIE8a6Tj19dp07jiVuE80Jl7QvAQj8ZKAdQ7Hj3hUQs88ruGMTGEZUhAQjvAVsyk
UPe6BAsgPyl25shuAFEIKfNkNth/hwGEOdrXEZ9mNdLQ8pu1qAMRnbV7YLbSS6fw
ZQ9UDReNoRLNLnqtnHcxymBRgma29Vq+JcR0HxouQKQ3MDrpBcyDp9vmYSHT59tk
5C9TlUo8ib7stEe5Wsuy6hF1vv7oCzanGXc8jiNfPrqv5FdvsPwhL8x35MZFgYgN
IbCirXwz+8tjqVRLglsgGTeym1JpOp4xNWAaXDvt2IZXqTnF+0EGgHHmMJ9bzd0j
ywS7j/MhCSDskp3vzDtW0UW4aulS0Hzaz2MfHae7iPVVJfHUA+0JfvBsbk0lXaFx
jLoG8i0FZzHm2jVc3uM119JV/XxAYTD3k7nYKKusU68zGP/Tf+GP9479mIo6o+Ik
B4jbmxW5pmDoFZcPELm05JYa2AnJPcBi9/Ti21xUM6z2FGz3KFX7D5R/l8rUCos3
Vxiitvncpv6ROLNyKSnWa2yE76iPbu4Hz6P9ce2+cwtmvy3b4g9jsc96PgF7yP68
p4xOfRFiIOki/JlC03QC6k0hi/epV662okq6yPnibswYV3a/1SdKNYfxj33xgvm1
viQaSptg8npvp2+G4bFrG5VJhAAu0pWQclMC4dC7Z7CCVP0tN3ZUwO5XlxzUpIZR
Xb3bsHjiTFmm5eqAlXjuuFPSAwHSBeaOS1guaeFyQytGpYEUeT3XIUg5ESffYcpR
IxMD39pRkF66uY3D43QgItT977gcWy99v8zlR+b53CJ9QyedBmjoVzEqylYebTku
HSM9Z73ZDyLt6xLOs4Up36V/CD5ODy5FPlxiHaSbB1y7XkoOonyhkV3LXR6k9IpX
ZTwDjoFxgPgeSh58iFS59IK14Wov+ZyvD0s6vUZi3aJWwPs823mrskT2/Pa2ryPJ
aX71k/0o/7CdfT333VTi6DUEm/2z6avndNw+du8juSL076aF7e96wT/8GfB+RS1v
Q5bg4qKgtmVloWjVvsrhzJCRoyTxVJLKpDi/h+w9W1PRhg5jaB/pxsxVABTIdOkU
FmtMz6ctuCoJ9VF8t73daz5bMGIhRNlEGhwojF9B5c8bgbsIBMA3hP/6QS3Iop/U
NNdNE7YXr82GvRdyUWjfOMxkJ1aV2S3pf2DBz3Np2SE0tJhlCz4s6X5qBBeY84dy
uroI7ySwVCWLnUVH+hbytmW5gsv3EDspLOtlJW7sPa+brjaJZ56w0Jsv3WvmbjVM
avijvNEwDCD9tpMaXGc03VcoVFH/93od1J5tFEWcountiNbCpR1js8JT28IEexWh
dRkLNGNDKal1tDdwaic5ESm577vAVAvjJVx3X1DGHNObNgSajWhuAIeld+k62fA6
hptVtLZnaubVxh7+oRZMQYOoKii4vJmbDLHipqXeS0nmydF5eFtgkwfdq8WoZ4Ja
FL5Dto7/de7KrGxDsuF3iHRFBXhUP8960Y4VOGZp5U1C0gVIqN5Hsvl/EM9Xr//8
Gg7tT4P8bzaYc4jfSlMD2zpZTlZK0p7bfCTIQWQbKymagXlJOFmYagulkuTKHPHA
O0GMTm9MB8iFe5z3W7k2FiDK/HEJ4R+7WeyGYJZslvRXli5KRZLTQP92GjvVvWS/
VLIAwLSgMaVQYJkovMe4QYH4pkrnHVR7hK23Aj+30SbbD7DYLu9QhX/Le+SlyQQ8
quY7N8/algDDDNaRQ/dsPn/FQ1IIAp3XHK/SOwIaz+SbFUAmo18F0CJmGE9SfW4l
OL2oU7qGlHWR2HPEgFGxYkdxSChrAXSQXlfjiBUkbQq9L11n/yFgvYOtaMUYpCfF
SSZFhM1qlYRQXdUPg3oWoR7F5zWj28iGl7GubXulE2s1w3P1pv/pahFHMlsNgYbb
CyaVh+vh62BaVn0oVhnVSckWhZe6XGw0awtEtW1WNd9rYQR3tTNyB4h1aiP6oj6I
fjSAJLROv9RMGSRTC1vlhnlzh0BKu+zZ1X8yUlhp6KnpOGJ+kVM7uHP+iqyd/O0t
LlwebXubmSDjNWQp9AF5CkDc1IaUCq5+/D9FsrFu7mbsQFpTJyT3kxk0Ljy/9h54
LYjvD8huFnav2kBwmrHvTZ7NEm2iI6RsfWHQ6kk5cffhPleQGj1cWCtj/0eQcuyk
XxYjSGm2GCXbXremBdueT2Kvt5HM2sxL9D5K4lGtcpPYj5i2YuZKAohtobTiPKPS
TueVKrno/yq8Ro2K6Io+tvxH5g2UFtrjOZ4p2x6GSaCkK1sELRLSp2pG4CjDu1PE
7v0ONOFWWicrZaYaH4sH7NjaisAFalwL6YDp6jwNSXPVdTiAr6RnE7KeRpPANneO
HhGviaq2jZwtH2Yk1l5T6yC6aQCOYSZBvYLvvpq73hv9JhxkeH3Cpqr/7S9XnkTD
WlJNF5/FTAC6BMrSFr8KfQ7tpZfl0OosfUDhqQ3H8g7jVBjv+/Z9PdU+yQmwtv99
QzDgNbnvCJNcy5Su4Mv1Zd+NdQ1XnoCtZlI//bvVEMHkc32QcZvUq7+ygmKRZqB0
cKCzdyo/PiZH8PatPl/o6nksROhE2NXQ42AlV7su0HODHpZbkZ8xE2bN8/SxlJWz
nRYpvMJCE3kMMHvkuIzQZYuj8jW1121IYS1EnG2y6KJGlB8qGu9+CPE1Ma9f1PK3
sR3GU66P5mj92PuJ0FCNJtvCcx4JeuXBQ0z8e0C3KrBSDSXGuSGbm9ZZUxupaxNa
eGzg++AyEayh0jp/y6m+O8t75fNY2tOAnaUhKOF7VJ/xX6cN1TV9jMNEzJUDqNpG
nAaN0OHiLm4VrQF306b/RoyWb/9AQBADn9uXqMnC4HFngrS5wop8BKekN+iLMv3w
pwoFtKh2T/csbFwTbU4Vt8y72TFUNVF7XAv/qMSPf6k0bBtV6gJ7to3ETOYYMpL+
XJ3BZeNb7oQiClRZrIJSeo4jdEiEMGt3Bb5c16YwAgrj3e6wAKwOqdHDAjx4O2SL
TZz0RzWd1cmSnHcSIRUyMThteonOf1/J3XCEb2srSfCCEYbeAqZ8Nhx0Z1iHimLA
aIpn5yV7gWgaX/ewMsuguEHLR3fOmUX/Oi9B3vTgunosCUEd1t0zDvrfwr8Aoxhw
L+05Lhaz3GRL/lFt6LKoVe3TZxf6Wx/gy6RgO8mN1+ikzkJvgeR1u/NNYxQzB5Pk
ajL342I19GQa7FEkbA924DOzG/WKYOwqicdfBlM1uqEcIuCCMVWwXQitqSahW4Aq
qNX6z5Dk6ObKapoZ0Wy7qvA4Y9wDx2x/AKWbDVHTj3z2Y3/gW7469B1giPlzYqAn
Hm2Xa+V5DlaKKmYm7I9RfDrrae9oXTK6NouJkFnhWrxosw+SpnIeAauYyRODJtWZ
evk1KJFKa/rg0tBHEbLoUjPu5rxi3zn+THhxFY70AnPF5nvkBGebYA8i2VWfc/52
YctEN4Q7sNJOxufYgweclFQediGt+GD45IpAIDZKPJD63LICgX6fROuFi/W2PKjR
ZDJmvAiSqXSo7arIplR0jEE6N/dmr1XV8f2KVtSXt8q60+HjrWACp+9Vo7Zolc1X
Z7CLzAqzQlHbS3wn+JruClt8YnfSnq8GrIE4+mner7Izh65Pl+8Cc7slu1xf9RF/
oLqhEH9XJ1Y87SsIZXenI35sguKyZA+Zgo6aJtjS/j88lTTSjPI/ipmtOoyB9y99
iBXagKRyMpciLx4YLfulgTerszDIFwdQlYvsyhD05YHTwLITVeEHkgeKw9dF+V2r
PInAGhkSDWWnsme4IYhyjTPinMkqfNkUHvoUDwT81fVjDDj0jBZitsiXW3uUVEqw
ICib8woDVtL9jArfiBsw0ldmACneC82UwgzK5CBKCqkCRn+Lk8q3RXhAU9KMOLWQ
3wr/B+DskAAFwgyZIaN5Bw/cznHJYnPDMEUQadjShu+JWx+kq/Y85WgkuJ3ohA4a
Zi1E40dhfDNHjx/clh/PEibFVHFNxW9/halyH7iJ7/wzgVupEz/EOX/Z/QUq1TXM
NQryVf+etcQHeAHVDUrGJrMDKHX6gJE7VezHlsftfQ3owAvWzU15h7Y7uQPnS2vU
aWtHn32/c6ecZdGTQkH9MWUR3Ru0KH8F4LXqa8GGgKwenEplh2jt5Dq+MtFcDBvC
H9TuP5WESh2ZMnffDcwkb/ON908LHAvlE2lJz2XZHENdEURy1iqJvUetTJMOqy3H
OAaUNdQ2Cbqt7LQu8DJ54RmBli9nX7JIFap9XeXiFyb9OdwXIAb8VObv/aetjod1
3/aM5A6NYb1Ywi8rzT/KHSRgYl8j8DvHIz2NOo5D41m3rk683f5amwlOkuP/aZ95
MeaoU3Oq1liDXD1JPxd80BCYJxpkjm8QJZAETK1GMGjNzJ4EAz5q3su2Se6QjHL6
HecXBZIeACWsVkXiq7iBlopPMGnaEsbB7SqEZRr1UtiavisGKMYVaKAeLiVfpnsZ
gkPNnoF/k3ZELCwm2tDCqnnESLAF3ShytnpSWsUcc83J+UlycFkqNSbgT+vgD3+h
5Kj8s5K6deVeUICSf6ndv7rpSGoc1szqySWAW2P2YcN5CTjz2pM5fZWrrllvvoIq
IRYCAUjEToRT9MIN5Fsm2ju64zN8eqyX/Li5bZ2qhc5eYNrBfHVcaY0XRi277Tuj
Y85MCwRHuN9JCtayT+WkOQlBoTTYL0LiAfFnMoXLsXmuUrDjXv8qChzOfv6brODl
cLxKqT0+0HK6GnisZiVJ/SF+wMXNO3ai/Gskug4dpOqSFJUmdk2yhJgjZq6chLWN
3tJ6pQ0DTFiU76cytSNXrYYzuq2nl3dI3UH8DXDKLdzxTaaA8Qj/pKTl1lgcePUR
DF3oIFycy/i8x4z1k+/x2xH0p7Yis3J5q5cBxR3SJRuczIKb9tGpwp3ZKQI+g5du
kIAJXwxNY95H8famjx6n9cEDgw6aHFSKZ20M67BwjyExKb+sz9nAaDNOReQ73JzC
g4EHyMbZ4GcPSwfez+ATmA3014j3XCFTcfCGE+TN73oHQZSuXea6Tm6Tg7WySOrf
fMehWj8JYdg10uSBW/OPrVrJ8qxUcBqPK0RjshvSg/XCSiGmNeXSPlUv3RQjlAu3
HlOGw+p+Aqpjo3mgJvVCg/ByUad/bORlKIMLeilaWoiQGmFqwXjwxyuQm4X3xQNo
9mejXRWD32nFGHPd1XwqGIMI/2QhVdv2qdxfFJQfGR7CrHOZWUqY/6bl1rV487T2
mj/ZKb9A9QJBg9LrbOAsatp8UZFIabuC4GuKVNeDKZdKbhI0qXlE/mwHsjdrlPpX
xbpMSqPmpezXub4D8XRUnjcyS2VXuVnuxjUs1/byCsjeSM1M6+aYTBV4THoJW8g/
fJcssWRu0VSXA1BDysO99j59EST1BF7FfW2i4033i07cwSGynUNSVuj2fIOUmEW2
QIczOa5sJ83m+C3c5E82DE3FE9hTkQW3AtKp3Z0QxnmhSE1QaCFaoI4v8r16/OOh
rzpqNjaEyX22NYNYMpWTUxFRzcJB6Qa3X2N4YDrgQZ9h5t+vTVxChr/r0G8Heamu
qTPDVOS8Z6efoY63SeefeLuaxXslHH6817Sa6jIBXfYK3MVWAYXlwz07LvMltmXp
bhQDCyxdjhG6F33wrgzB5xCTFOfV4WzHnmGpWHti3xaWBap/IdsIMiSz1cw537rP
mPzrkLsA3QOEoUT88uBIlKZkqe+zQ8HrpsyIJ6F1DOIRRy7CXCw1ABhq46iGZXcc
tkip24+P/wmklbS9CStCjftkcbTU1flq9BuSVzOgPBEzLHYQoP5mpbRpbWjDF2YG
ALU45f56HUr5svfLRwY01PAIpfAho1bvKB5mFRclt6vPY/GPFVu2ZgJOxh1Dl2el
fH7N+8i0B+NH7iW7OguoM+0+nAEJ6Ti7LUR0/eolgh7577u6K4F6y+ovfq6SsuLH
owlsMz6WdyQYiLKrxggjhLYNqf13QwYfqkxskk/OeucYQomekPMq/ZU6bScUfxHy
LGjxqH3dqhjIOyHv1Yk8bR/ql7tl3psr6YEURQclHPs7epXALp0XlwhGDN8GCRXL
HBH2v2Bi2aUxggHDr99Dy1jpxMroBsvp0GY1P0x2S4XPSMFOJkbRYHxgCfC2fnj+
i8rgfAZw9ruGRsWiPqmeUWcWUsCle1iV46Aoqr+GfKjER5W9rf+MACPkckrRNKiH
VX4LJ80yxTM05xPTo3Hcvu0nptb3mTyktBNzOXXy3d32tXtYDJ1BsWfz70eOe6RR
yr1pTFsHpGgOVhdvsFTRauu39HP8tNVMyZpIV+w0KkW+0n4eoQ6EMMMtEvNl+lUh
HIwgXnv3H3yz+FqpRm1yqu/p9sJU4sbiAgl7BqofA0nLWa3vRnxCqq6+Uu37leJH
/4U5k2siHP9tmSlJO05pErIePPiJVANAYepeuVdjl5bXdY5/iXM2vbHpPHCThSRp
yc7KVhcnf1kMiuKIsooagOht4/W2r3pI/I9+B+SA/aUpDUmt2xy11aSNLNGfZD9c
LCYS8jeUjZfnvq8w16zYQ5yzPXhZTsbZh5BGqY12G5DYI9dBBoAu/23lupD21l5B
NoYcJ+3K16HbZBsXV6US/p7CypABWSXUwHuFSO1mhq04+Ig7e5qyBJM+oeLPjs3Z
8YWprGr1dp0ghnfSBqMgdFN7OxN2H/1iNYReRqdBzrrF2JZBXZEt7kgIfhtUes9U
YC+gGQhJZUg0TzkMO/mNrPzNYyZSklqlhfYmsdvvzzI4ojZOomtKYa51JlGFhvfC
7YnxhTKouwer0P5m3dplk434dPhXkWBuZjug3PdsYV8WazPeqW1rdb3EW5TaT0zH
JZh4+KDvZdwZR2QAmfx0iLsdtCoFhuypc1S+a9wTqdFg7cDsY5fcY1mKT4Zd+8Oe
8S2tEmWY2Djr2SzHMcbsLNABfuvsrQgnmr/cyWhoSVls8o1blWlUBtv32nCrY32D
R2bxnhQ5G66zTv/sYapAnxkNRHlh1Y0vFucbbUu6Csq2Mg+kOHacmxh2ISzuohY9
4Lt1/5dMEqwsd0e4CrbprPpKk+n5MdPPQiJXZXgUGo9saQ34K+cTzOpB5dWmuwdk
uht+UxjlvUEa3bDPY0Jy45EEHo4LwKAW2fomNIKAN7pcVsGOWp4KXKEk7+kpVsHu
i5OgpFjSevLe/wDRagA1g4rBSPFYf3qvmdSa+FB2KBpegl6oNBrYLMCeOL6tIGP/
RwczZFntD3hKczpAJBsz5/ehvpeK4sOszRVAiXeI93y17JVZc/iIadSlk37ilRM5
qClaYeiybkSEoKD7BMLJ2PjWyxuCHPzldXwg6tKGzmqhhqjpLFr0IpEVt4oc81Du
TwuXJR6X8g0XuFH/Jkiu8fptHY/uKCe2U++kd1fdvHfC35UFuMaBZP+gtZCmhmeM
ZuQ0LaKKzn8Ly1WaEB3TGjefhc2Z8ZnMNrdKUQZHRlbgICGOPWG32bSCiceH+m4w
yXzAEWrOEFJOcefILv3nq6VFfuZsYprIl6q8BXWjtG6gOD2hnbEcqfpug2vfAngn
bC6bqQk556BdWQ7izSfRAhlGNYGYxnKLSiaXKXq3zxAXMVp4IyHgM4wx7qcH9pGv
gbh+UOE3Uvuc6mARjIDCIdpSdo+oJSj5quqyayzuqlDIqJ0jzr+FVO8kqhObji/e
ZZq18TzFQ7mCUNIerz3Ml6c6vCoJwB7zdBkGGGJzublduKLNjY02iT+n5DjMVsLZ
y0uqRjasIzPZcGk6Dan+m/OZwSzrGvaFdYWmBj/TA7DhRwfKpqNAKjzhDWXulMn9
U5ZSm6JM42ECczqnTNZId+UIyEBJhgiSe2rQkFgKUwuLzKuSZtPyo1Ove61asgMK
oUwGLWv1W+YjS4wdeViFR/UHhwZ53+6cPdVumRXSVchX1cvVTuA+NweAWcczzHKa
JTqfzW8JGEjUjvLR33t0ihNIeO8S2jlVFEdR5FrKI4ZJ4xwWLDBQgIhkAsGFiSs8
KfizuJ2NzB7DgcP/1oWi+ExdtgdoG679PjM48rPn4Ef+/4RyEiKDLV5nZSkxC5+3
xHipkjOy2lXpSBFhSDov01YLP3f6ZSrDYtiGoO0HjpG1UwzUAjjRAI68CM7irfcY
CPU7xca6osAbz6s2pUAjWHkCR5Rt46+8fz9lJPnVVtPbfHVRLElEsYF7/LFkn7qA
lrwvtJKYw1O6L4+3gsNWffQRr7XOKfG4BL0XdOMFmjZ1AiL3Q99bxQ/DpYTj+LCD
S8TTdlcHGiP8xZKkjMDvknhmJZDemspefp45Iu3XIfGlE9utUbKFRudyCDg2I+WV
GvkzEKQRmZ3USp+2oNZrm9Kgzca2W9C5hHo27EhOdp0SbaLln24JmEj+zkAXWtsv
HwVdCUnZJho2nr3praziQyMhuBH6nsDcTlqW4C9MgnBDX8sOFsvStUvthInr9mYD
x/dWolUYZrMN1K/VxXKFfo1c64fuVXlYT0G7BsrgoQeB5vNgIfzoFkr4T50D1Ayw
1EQlPMdE7TwTHj0YiJB4gdU54n4dgOXr8UvIUuECJ8gX0SiRTa2Nx7Kx+DDfMML3
iw/VBIbKASSLRn9qwhZZEK4CX/1e3+l/kbrFrCFilyRHbIdIxET22FpKjk5AfGhL
Q0AWS/lO0ULSxEdVPHvVvza94m/R0xdpK4/mSDetfdWh87GWOsNk0hW609DPp/ie
Stz0t2MkyM65o0rkalaZA0PQy3TtjCfGHQvSxqvoGecggMbnk3J56AizdfA1LuY+
JJW6Shn87sUO36brX0llTw9KRmGf6Xqizs2oUaVu5laQpILVskqO7gLT2H0RmEt6
YHkZcGa/O/HLLm94amQOjxEWLJclLjkS1C8UVTGM+G+yQrHfJDW84SKUCff/Fz6f
Rza2BwftDvVL6x+nWXbeAb72Nst7f8shPn9NN5mYBmzdEeHRy91a45VBAVBtBkn5
vx2ZPsm5UUWUhZigrH0wrJuN+6MBjv/ADK37CSnHtwi48SE2XwuqUeFCa4vmBEl9
WRVCES6IRpBkVGGCveAF8omUTzD8Va6lfgkz7FSJflvZsor84zYvL/R754jnOahw
qfj63WBa74KlXPnP+6qVvj5+/jBzveR8y9Xdbb/daU/lFcCgUCeuEFzzYSfJ7sXw
Xojw5IJbZGZKZNzH0zZfsuCksJCE8l0QvgjJdIUd3fp9tqUlreoskH+kD5b9cz5Y
Ir28ceRmd9NA8vQclhRevO4Jup784Rje0+jikyDbIlYmrOBTqZLTc9dMZHEdOsyu
A2e/madGleL1BtcGdCo0P2d7YR/wo4tNBWFaA/mvcBERWxBpsTPBUEzR0GusPJMi
MtrAHuUsjoLguAoXnkw+vXzhdeO5cdFQ+9Oid1UPfT7AEV/JuW5DcQKNjlZLVKYe
ssDB5EP8YgtI/BttlM+RVkLqU/urB5MaRJz6J4z6VX9kABmkgLMP0vGx8Oym0uEK
deDFYYsi/vmMhSt1tuB9aBxOXxQzpRqhbwUQHSE3ZE1TOXHDeeSxlZK8ZGR64SW4
4yr7Vox8neE+QpbZ2LHR9ehE4dy72ZQEZMfVvAxqvPAU6g2WlM0A3YcamYcbCfBk
Wm+VuiIIgld8mhAEQDph13AgB+TT0mkq+Z/ofq3pJIJ23HQHUyElTxTTAUdP5mAM
MzcNbGNoQtU48shrJuLNMhyEuBl9r3TulMNoNycT/zrr/7mOtmC8GD+AJPX/dwpY
pK0Brw5Zp/1HE/SP9FHfXX1QwinIYH200bUy7vVo9w8Rpraii7WKEW7Jaj3fDKGS
UFl6Jimx6beCKJXosOvdSKmADJQZhD2GENMfd+FEmLxO1DREce7QKnXbu9UNpFoZ
mJDEo7JxAzkOQeN4ipHB/nYq+MZ5KkZnkZMiqUaX546IeSbH1/BfYg2bh0WQmFjF
CCeUI9Vqyx9p35+5ujdbzfzSe+PJP+zewuDQNpGpK7UwBpTy3JWqqfox3p2ZZLcA
gG4yxdBkgu5zz7DdOE0+x1SIGPZ1FIim5uCrRD47vHE8wZpM+yLdX7icQWM4XcsJ
NabkbBs6AvMKzNTcuO3Oxdj4UFCCZUWtC0KTmUNNxBw0613QrLQ+8vzRU0pS6NcA
52Sm7Mig4/l03fE61SF797sVsZoIgN5YYu0vxLe728B+wm33vM8ixj7AArlf6+M7
1UVtr7is1sw1/NgTczW/lkpis4b2/MxLwyeWo9Y2Cgnuz218dRz46XC5ZAuwPD1Y
SRy2BOQSrEjVaRqX8lIB5fK2ufGMZj3aYGH514HcPxSodjyVnzwx4AqykzPpK/MH
/eC7TlSilQUg7ateI99RePvpMKnVtftiaVMJQs1+592su0gTw+QSaZFRcy5zC5+S
cR9cmBxwBlNBgMLfHDGHXcE77wU3PGNWWYdFFD+rwWaW4prBCOY4pZ+G1U/OYuID
O/1yDb7wDYhRDJcRk0RRt+FoomJgwzx1NzuI6LOVaT7q9aoLZgNGP4yobWBEBTbM
LXb5jDbf+a10DKXNIxhQKjWeC/7VP6OIhIKJIKyE2ScQwWJ+6y4Jzd09Q4WQnKKm
ugsJfQBt+DOlDnIpq1m0mGSOgH1ZDS5qA1h2OyA+7dFVKf9+lTeI607/lGB55pAI
NsDaD4O/hpyWVdrNY60TDEEq7zlihNLCoWKzI95hCGabjVZ4UIcSKixgdJ9ojUPy
zPeLh2SPc+PrXGh504MZFZK0yeJdXF+ZHZgJIwVJayhvQZy5yK0dPEvyIcM8MHRC
FtPGo7ylA+yzoYa0BbJOr5a4Q6X0bqwS3eS585Tt0cv2wWRP6iG/mL+D3ZQI34f9
7zg6hkCBTteE5DBP9zT8dSp9InNKqjZtlFe6FP1UlaR7YN1SOTZuAm0TWhjrj7eS
1QynGxf5T56WO8bUjZnkwB3fJY4Pq+DT1FbEaZWVQIv46y41ztsC0MG096mNZS3W
eFkjbA9Fgh7wVsR6dXptrPcXn7k5mkM9vv4meOQ5DDjpzieWle9ArBOMoeQCn7z9
nu+9Kr7Yc0kfk4cL4UwqMr0djrzMvwgwKxLpuaF/8XePksOu5wVAMgxdQUmIjjJD
cef2kccx7tfVP9QHhatV3ionubQmU956LzoQg2dwj9ibn8JbK7iKMWkv1K99UnHt
1PsEkxA9vCdI+9WQtOoEFnTWClGao/X8EDul/uud1huNnmJQvkycb9N0XeFAhtT0
uOGNZk1tksWcZXNWomTrpdT3/xPLteimM+72GgsiS0slaxTMfZ1ze43ZmkNHHPy2
uPbWJNkf2AOfjI+4aOpeD6GNxPhUVh6eL3gpQDp7As2kyY0tqtgh5UfUYUNXwV6/
EtDkezh8PeC1kJdQGzH1qvD+c0yDM1Rb4mTO18WNQYRmLEitB+pXqr7zF2xlvzOE
8sx0eOY1iCluatr7JYD8nfLzgdmk5h/mZWXDAqnM6v2IUqdC8JFyaUzRlD44ACJH
Gmu6m8+F4JIQXVIi0+Synd2XyYtYq6hqx4HhHRDehD+9ctf84R4lIR4YiT0S/PMF
7WY5GZLxdpQOjO6vtjl/PS/pn20zxor5yUwumCGG4d8do6A4dfws3Nh/sseK74qH
yBcF/U1znAeQkHCYKLi3pZ/V+Sbq43Lz8bireZB8rHUao7m4K9zquEWs+OI3S3QZ
e0C3fPcuWLXzhSGvxaP0XNzXlhi2dsKwGmeWcdBv0GfvtHhMefUgvkXEoZbWlKMa
d70GyS8kfDvM4ASbX0kxE0U2YFxXkUKY0sVmILHn+n906I/uZiC4BSDQYKlJ4DAU
LcRlB3do94fBF/auLd0Sb7IYwbq8gmEItkpE9c7BDGPNXvXp1Zg5uY6SOR35LnrE
mwwP5Ux+siYLnvDq8d52ggG4rToNBwNABh3tfD35CbqaTmV4OkzBzZzLnnpUxnKj
QdZgfrfdV7MxbiJS+ndfdvL0zpBZ9NMELMOM/DuCoMbuYo2IlO4FjIGl9/VHkJyk
0cTTmwUd6VQmJHmDjjcsAVFoiMk2ptqxL0xKT6NtV71J+23lZUlosUoXDYmVEzVE
uKmaVnhOPkSImKDkzFw1ys3RNv9QwRtKMwPWSGrkLURSzV1yqIxNuQJJKPvO0apZ
1YZjWpYz7v2F5pX1ToVoBUxvKOePzNnHNopQYwhgSRNkKyrU1zYG0oJUGWWnkeiv
9WhjbLLGOQDrwbLlGOzNfG/A0Be1YuBLqMETTzijYBw7EV2xiIw4gILP4A9vHyhP
yopyxUF135DlQlALmTI7K6+aC8LOcbbvWmbyUcvvsCzaQKiEx14ZuBxWykkIpod1
WYlH5OuIWxcfy3ux0pArKg7WDepJLCd5TDw+ttqgbyaISjyGDoZ8zRJampAglx+4
vq4qwY+eojRtWKRjXLkqPsCWCJLBnYRJq39w1/i+VEA5q5FZJ6F5UlE/+MhmRwpS
/X65eiDeQE/JT8NgZfgV2Z9hsgK4k3TBtQmo/HN5dx7QSQ8Gd3cYfOHBWCkDZMOW
nAWYLQcI0yAlACbmFNoNR8Z7F9bhzrSSnsuYivBvYL/Qda8M7lpYWjLDrshYgyAW
BiFIDhbmQgneiqd/Lai+QrzFFBnFDBQ85iSBYKSjj6I413adD0BELML+ZrrA4Ccz
JLxXyfH/a2ULvgjkxWUpFNhOp7+LE73bEskgzEX5Xkp3CSfbb6/FClRYIRZPz0xY
zcakrvE7JZXhd3/AkwuXAHieQj0iqX1BLf61j/LssH13x/E2/s4Mo60tp2vtzmQI
5zwvmF0tJVqUx9SPjLMsAioYP5WCWTAdi43ejR8874vpeNyipAxHTMxYC/+wZ1tF
0m2LtJ957KNEC/FsglGb0BWBZOHBfxUe0Zf99zpCgNkWa+yuJsbjvEgYUZBy97uJ
Xzmjq9MCxq10StznTd+hAHWlWi4MGv0lHgBYhZUiHqwjy0Wt4uHWTt9hJKIfRxjm
Sl/6pdzFJ67dYim/m7DyWwO2HS59DhrTXuwTk1PVZJ4DAXian94dsrf/xqmNyyXY
R2bMwh+MPBvPoDX2Qi3eiVPpccl8e1KKXmVgbRoyqxpK+7VREQNal7zP8OClv7iA
PyDmuUL9A5+VbF2wSKsx6Pntr1JJYkHoyl0eq5QhSjXogGGyQONaju75f/vwWRcM
o/rMgOVaTG3oIknnBF+uvnBwKEuPx9lqCCFwEfrx/Iz6Til1idZ+nnsjOziSSYt8
mytqCB5fQQMg/XqYRNtCcDNkFe7c2zjIEFfww1SCxSt93BFRsendohiKqsrJKKNz
3b6B/koenIb2cZTJIDRfh+uIKDd/iJFCSfz8UYBTI8g9diIeZKbwr6LkYmCF/p9z
Wyy0VSSqmZX/gBzuQKYoSvXOP3pyC4PL/XDLC8EAumgeg70xX+Kj49xcKpV0EXNV
gnh7KcvDaDbDHlgJTb8t+TileJZ2QYyiAz8kB/XOYYPAuEBsXlyY1zb2zu0TYLSh
pazxfGCYkq8ETLLTVCo2jEe+9GAPPIEcS21RQIAOeuswi1r7sSdUVzzW8pG1kn0i
Wx6Qq2bNkoZNqeuCk9IhLFxrFoSJciYq37gaT9PzQsqtmbEXtKKvKF7tGGk7VDvP
jVr4mYlMMX07cRCLiQQvkDVgq/IIBXny54q/X7IAQp1Myg/I7dbQZstwIqYgWGj3
tNYVGe0/IdLkaPXW2b4MPxPHoLK+Iy+drDfxPS8Fl3wXlosbOOdPpZz1JkZQB0Sx
ReY1X/PXWJlT+zCuyZrx+fEkdxvcgf7FstxHLDq876ukLbC3y3uEgo2l7WDCaQsX
HIkocClRmg3sn42d/TJgSabWObwdomdU9Ujnbb0c7zYxTap0iMujwNXHGGXBn9kw
sGwv97iP5IeDUvGffDiAYPvz1tjiGgKVVvEZzvrlSn8ZWyHZ54yJxKLGm+jqC19U
ujMUGIwPyJlnQMeoDt6SBcM9pIc0q8NISSbTTsvYVfSw8qXjRy+fhuKt/3ufm//n
ya4m+iMNoycby8iC51QpljJrxraoEPr6lUPuZZh/FD3n1lrGXbcj2Y1EPITjoyl0
qOll/jLVLX1FvxFCNOl1fwELqWHb+HthU1CQuTpwaDsrNiQzElrKqrZ3+J6XTXwq
PiGvR/jX68BodjfbsDqs8kL54LVtLBRG47y90mY7uKkti3X4JGQMhSWMfeQq0j5G
PSg6I1nDBDhjAk5MxvcWvSZcrVPndMtVvBAp0Bulm+Ue2LhDivlc/sFK9+tFjCw6
3Eh+4TeVY1Aqpbpvo7D2wPK3LY6gtrpaX2okuX5sExDzsmrnydw4/u+DAK8SAg50
ndLENxudGh2bgSXBbRt4BJcsqxFDXpT2L5TBz9VDfW5ChDYdMbNeBnZ2ejYgZF03
ZSwA/oEKW1H1lOVbKxMdu3+3QeXQnMkRCvTrYD9Kliwl8bu3Qkk2e/RC0deZGA0A
jbydYGb9wqJq5BsV8TTxM7Z4Z4yTYkemqa5AMX+BNQ09/CI65LS6d9Zsn7JxPoRX
0rVdL4JHBZI/vf8wAnHylbk+9OO+OB6x9cKs6mjAQ4cPPEoswY1TsWXn7N4n1Y74
t/HeYzSrwB7Q2V83Pmu1wbkZRdCcW7JhhVrdn0esssBo0zcqOxQZYcT26FKE2otS
nlyGpfBfnnPSYyqLPdBtCZVyS6JqxvjZ5abGrFFwrTUyOzffwLhJsYO0EZdfzMT2
fxXhRlUHnjvWTdVcneA0be+Ndz0BzxVnGnAbwciq1YM6sfHNdAP0YgciAJb1RItT
yWWFaqVDerywlyWuE9nDPciQ1vJXfoF1Mdgy4zgUR2EJXsfeD6/xiyVXeut3FATn
1zjo5N1ou5khmsqhJdslUdK7N0vIxVc/6Wx5pF+VOUIqTc5j32ydhpXffJiH80dg
9KAWOPh6D9ftYXWSqBZY1z46kTVIhmQM4D2IKrq/Jt9Mw8RnhPNhDvulNeyM0ZWj
QaR5P4vi2qXUIoOLD+MnXfOCOBPY1Q/f5DIRYdfcgy9v6T3gMwqMRBZ8sxC6GXls
tXh7zNp/HTTErEwr6HyX2zW8kw8d7mwFTDDO75tmRb3bUactPHzyUEkbrzk7hCSj
/A1nikPKXA3jrL33gE+X9sGSTBRZ8tIhxi9EXuZ6M2LZ2iNu5ZmO/e32yG9VLGjl
7ZomtrtrONfAJQn7uGQwXkivk4TMYB8QNjh2ykiW+RbbUI+2NWmTt0DbpDGe01Kp
+Wq3isrSCFYNaKQ8PtsBOmQ/RKU++YSCAsTNKRwrnxpBdlWCxVcLCY3EMxr3SlAU
J4JKA2qEKzH7oFz2bHp1IM/ERm9jwEOc+i8RPqq5HprdQ9TAtw1iLSfIFcLPaX0d
O+2OUdviV3Zo8/yxciTdkHa/uXdsghw7XnHuRtAQlFyOI/VVqXOf5nLvJLuvI6mm
tm8VnGPneOb+IFSLuybFFbOvC+8TTcy8nwgkYoWG4oJzAzzH46K2ikwBkLqLma/p
jWptw410C2HvBo2xm2tUm37+dEBgs+qSNxRl3DFFe8abdxHFv7azm3obclBgqqmv
Vpagl4i59gApeS+Ve1pdqfU6ROP2722lLkmEytDX2FhDRJa6GnaFhyhvZ6a3bC66
W14EFqlSvXU1iG1PHMPzEPO/J40eTwKY2zlrBaQSqOxUI4IfZG1od2G1Jx5pSj4n
fcGiD3ZT10xPi9wXGc9FdH9Kldyv2NHklTibABFLC/gV/l8s1PkbGhKn1EqgrSo0
IV6bt0DxXY/X9NEJ7nUUT3CTX2DwvoyI2eX77RGdWd+FODiBmUutJV4lIDcabP5l
LMjiCKnxDWh0m4mAl8SDc2/RahW5OyHDahBI2Hrw5iKfecDeu4eJ4yISg3fzgZsj
7KHcDX4OmlO7EQRS6uJwr0pBBiSei8Ys+jpVWCHUhpwEYGIYjriiwUL+C+c8Db75
B89HW0d5FR6SPwLUg5bP6QgyO1dy19xXj3OrshXSp7FwCjTp7TYyD3Cs6iWYFrx2
mPNOYjdwT4pmZiJ3exsrL7cWqpc3gBpTRIEz0Uca5EYmxVelZlgya6d/nmlpfEZv
bNeL0tC9cdL/XcIPSTen1pg/pS8xOS6339fIxy5cO/In74Bx0CkFba+kbFuP2Kub
tOfbFR5JQ1WJ07DhINpJyYDOCzK1/Ot7Pe+FJ7+qNMEPm0N6OGV1Wvn2rsJdclXF
AmM6YQdIxYAysgFEpUO+rAtTrWG7mf7/0mZ3sC+kfRBU91dDfRmxyoJyO60D1wVg
BAg9g0vETl1LdmVLt54nD11AyYdtrYSU4gRwirVZ/Ub3yCUwu1D0NnIXtJoesYsm
bnBJuwOMsSVs8/dwf3IeaW2lLbO9IXFVax12G9+dAswsVQnnR1KcSsBU/qxyk7Ul
8tHatl1lCesUSoUqekxI3HBcvwCFxrypCgHkvisJHvA3yJyJ21+CihPXswodKWfF
KlduZccRD2U8QRdYw4x+G4vP1ZvHvRZNMUSnZ7fwWJSyyhh9YFi3gR4FDH719nY6
31Z+xf9cJLCU1XIduH9F+COo+Y+oQ1xvTT4cevowakuHOQLXBRS2AcrZ2zLKYOpp
x19LuxK5EAUtBpSzpX5R6/FHcAZ4iyzm/cxoYJwWtrACc5dC1YN/Jsf2PVyEm1C1
f9LNp5LDbiOKFT2jT6vgZ/ruro3DfjZzVlAWVnH2S/ubByA1uHnkUgKIBsJFN/d8
H+XbOLo080G299namZfkgimQEDfKEEkdQFlXDCeJEKFZPJ6JzkePc7iZtmxJdBGe
fAncqvnjm1FK+xiS6XsRQz8LvPzAKCDqu0m9CSXD9vS7OlRVIuRE5RUxchjAVlXx
1MyA5XFgo1NicX2QnHa9T47ElYaBlDVhnBuSRz1I/yiolYP3flu+4UpNs/K6Pivc
tpLsNCERYy7Ah/QJxA641gTeJWXme08xbuxaQs1if+9f2R0pcP6MaWAmAu21lXqO
DqO2p2VtOqpng2xEmH0qjKukZOCewl9qVu0xa7Ht1tPer1/NkwzsvrF5Ym6UPxMM
sAKT54xe4uwSIQQ14rRyDhejBwHAAug7NdKSNuELK6jf2YxBaXYZ4+T0x/JRc6yr
tqKGE0tnhvIe/lo/UHOdek5lAfHnTYEkesPimR+kRUVbH2oW+FY06qK8bjZXJUoh
ecsjSTiENJBe4yWdtP4sh3B4lAMXIcZsuAlSCtsOioYC24exj+92en2cKrVoDxsS
vJMp0TUJmblyZ3wjiWJujhgWuBNca1Cd/vRUSEl7Sqh+GjMzQM5j2oonMHqs/VoE
eoppKg9W3iZo6XX5W4ewih/GwpJkzPGxc/YMSVCzXZmga3vQ1FasSaTddx9VzyBo
sW00CQAnBZIXjfV3mXpf3x6rztNYk25+e5cbObxxxMc9kcrBhdQ5Z6EzRqIWquBb
KPhyk7ZJzbOb+8A/cTRtwjNtUbuEL4b5v9Daag4aKTDTj3lmT6uuKZfGhz3FRkbd
VXXY6KmBFdVtsWYspJa10ISEh/0yEtAF1rLvMAyAHQ5/NNbGdZC8U1kBqTbZpJ3f
PTB1JjpLyAtaCh2ZC7UnyAejdbxGgp0tECzfwcWzimXLxlSaZKSKwcGvBIxBJz9X
a7CY8JZbWeRgOWapg1c/AnDpW0hhCSAa1IvyaJdbyNeSxxaMFJ2rVFdnsKD5OZ95
QXMt095Vlo65bgb1TuccMwBsND/H68joM4gQJFV5KwnWOYvYs6xXfRqyjUr1341w
33BLmg9+aMKqIO74yakGkx0Jm7uPwahVy/CofSaeLviLVpbZXCCXUW7Is+Le5Yja
ZGhLVBAYSSlQ3GLV4kzkAN9WFm7KznVg3ntdKczOkzAzoWI1kFgLv4nOH+ybRKNx
eyZfIfvKU50SVuN0xiLToTeO93F9TQekVQ+86f+xTj7pY+SdAeeucCeh0s5icXyi
bwvLi7G3MvUQAsYvq6h2zyP7iNhHBP6IVE66C/zoGmnNw5PgCHG5/S+dhqz+q7RR
9hvJ463J1Vp/5QJe7m7OzuBmiKiGtxmNf9QNMGZvi3dvVte72eUs2scAV6CRqYS3
1tI129Vn8y0KdFmGsz0qr+//ekxneXBcHswMo4mdOeAL1/74eXmBy+2gDKZyIoXi
/ZGTuIoSn96i0jgQiNFzQlVcTrcJZnzTJ7bcC+7aIZItfuOCW4vOdNkNeF9oh1j6
wYpcHHXyRX83dqEl0LtDW+dkFLpo8O7HAtr6IvINZz4SJlLmSK1Z5jD2qZXEkpVY
bIPrqlRiuTnVGG0ZvagKGx7G4l1f6KWZYCnq8kmHt7Efkq9KeN+t68sNs8lORt/+
y/L+cr0kn5ALMTaqTW/FaIL4warujfJw0KcXpP1/Z9I/R4JyLm7awWk/z6+I9zrf
Q44FCeTVIkhkfO08MiTwR46aOduQh8eMick9WIt3fYMQgCoyK1/n5xTtAfP2PGzt
LIuXI3pF2+/c/mGkqLgTIFuxQ0EVJ51gNd0GN7sz4aF79jeDJo/LNgCXq3J2cmog
phX06IJN+bAh4lru6y+1Yyd8iK2Z2YLxNhU7kWG8iNqd1YbO9h1IvTnmcZBVCRml
QNwpTnT8q66fjSyJn2tU6sJOxCx97BKgqVmNE2OrYcUN0CUgTc+Wj8KcCecdYDnV
uGxF3Zyh7j8xq/mP6SLJJE02OUIl3u2RvCMNqVFeCiOqjaNyEsLK4JM3vWr6p7sY
iIW2mFwHeviVNuvlTq/7CR8S/nXOcXW70Gs+bwDw8jHkcaLPisndVAg1OXnwIf7C
QKxj300fTtxHaGxzbB2onYWeB2SP7TJAFQHWAe6O50R9aispNaH1u0KKQwCZwI+T
aE5MH32xHgs04kOsl/5FCZUID6Buge60817IzJI6i78ExuHFxfocCJAJ8BW6jY/R
RazpUy3KKK5mSJcByhAiZVe8P3eG8FO3htLTfGCTutbcTdYgMlWyAhiOo+ohSEbP
L/6fu1bJjN2Rriverwmd+/1B01CAH0l+NJ+SIPihukHM9vmjynYPavMomIDqZ0Uv
dsUYesCUgw+iWgZLlyXDfINQm4nR2Qm6lEuZIJTc27q7hd9gBieWyygYp6FnXs/c
fv25Lpg0PFjFkBvgAXYAkIiJjW8J8/XdYy7I9d0uWCAejeo3YgGMhCZfl28hNujh
Ra2ZKjwX3L1EQoF8ZWdGslB/5z7VLXNtyOlRWDfDOKBAM/6sHDhV5Khp1p7AVzgE
VLHNx/z2Kzpt4cMXXCMkihhplfDjGTT/1nxtpMTP8C9wOYilAFyipZHFOZZXbh4W
VdJH+f7XFUU0OlpkvUBl6KcyaFjrFsZ6b1Jpm72Jc2bRBkHx/4Z+rZK8V1To50rU
mnVRxRKvYCXWUnGrEN99o+iXQ+pBIxenZudrB3YYmh2JmaDxFsIm0NB1IqJopgWP
Ih70STUGekZuSMaNyxrtHWiKjBgAcsAxroRFLCIz4uPoXJ6zhEEdYEkMLn+gUOmH
55heCXDFKQrYHW5is1A1On6IymoGdA7ZMI+CdwJmwfGB1qOHCBbWumPET4BE8bUQ
Zn012IUoSEbzb7vx7n1Wj7D4t6gOzRCXQVpGHPEIGIUSOi8lq0BaNwu50hvWnmhc
9XgXe7C5/jCv92XxP7dGVoT1oLzlGna1CvzDLlLM7rNQ0Xu80yUYEcinNHfTqhtT
HhVCzdMmZvwxI5sBgasv5fz7qZaINFpXj4SDof5dNf/fQ4OU/cc2af05aPqBuzEJ
p72qB9iQZKwEtxN5A1XnSd6BeXGRifvAJd9HyOtuBpaAvNGinEU5Fq/GzZhB856U
ViLwYGR5Ftkw/3j1tKxYp5DGiuizeJOsB3ETFYDm25VwHhbDmPa3nzzOpmHnr2xE
5EFSqGH9ZDRU9c6uHx+/e3BqTzG9ukfeqKjs8YbZbDCXsfZQq0GXKI7qEnapTVee
D2r0VPix3nMxsKCrExP8xV4+mnOalI1t4tIcI7Co/d7nJpsOtNNm3gicDY5WMLif
hbId7BdRuVb0M/SV84tJUQRKhBN3Rs2sYyvTCjKYz3mq6DWdzbqXb20e5Ib+3W/A
bmPgdwB+CfXSYdqzMf7f7YBvv2NSjc7zt/vybh3fQTJ531KQczeajayBIBVx1kJM
9nCKJpZmdq4uXHAIjG5t0wcRQ2XwKqeBTHWiqzkUt0NtGfG2Y0Tk0yfUoTYdxiAc
jB37fBIC2p9AiZIFE+tBqtrNj3Dz1Pl3V3TvcLO3Syhd4y1M3MKW/ufiGPwXHWne
4O2piRIdA7RkS7Th63XkjPd8iC3T8Y6man/UIzX1HpOi0m6r4RyEvmxmQFUH47x8
xmv3VIu7qikYWtutB6DBGc+IeoHV8hS5k77xu7OFfhK8qlOpVPvprWusj9K16AvD
o5fqfPKlrKVs+WfAk5/w3oUPOsuWXWk4bmZ/UeChCrWNznFJ41FUvGSVq0E/NmKF
453S1eCwd0otYVmn422FGmLLFf8pWG2UfQIVmqWRdcf/vve4YSfr7QkqK7ZTPKSj
i6i99jFGh2IKWVRNsby14BKJEFqd11gxPt8VSSrwE1aDLlfT1+wAYvlQbRq87xPE
GzNjr2MaZzYb8Iry0AUJ5cBoraQrLDdOTwcuTTpQXNbNbqo2a/bSzH/WGN/Nvuyt
R7Dt2gLNt5T56IKHDi5ulqI1ewhIn7J71akGCfWRcEajR8FYFpviePieHufobm98
T5wPXFfOyr2RBFenOY/w0ylJHGmdMr2IDEBs0naaOz21mjGvel/XsKCj1N7btSyK
+3Mn3UfpW3iWdMhUg5fQZYlrysqCgKe8sUeGQmjq69sF+ObN6Atw0XuYexNK/3O1
uGQTIII6OMvlNIv2AxBDL5yg7c43d+MgBUUSdC/huaytMZPEdCXlLdx1rkFM8U/O
yGufIRARnaEgfcrfOH7CxM9ydfFe4l2jvtIp1aq6Qn0BoMl03lqwsUWAe59uNosM
36AOolS5Vj3aKnIjFGuUbVIGriKWRqXWqGOAceS9MYnzmdliu/1zuHAaRyPSYmWI
nCQ6YPG4vOCoSGtTMbwAcDQCXmWnGx6WvCqs7j9czGt+u1V+ei3auPsILOLpcAFS
8rISJhmhrSN1n2SGHoAGYe4ykqHOc+Mp0YCtrqg2Bzy7Pd4MdcscMGpLwFi8i1s4
ALtBbyKehBcZZA7PvsQo2ov//mgjfNAPWCiyNyiyBj8T/b4i/vCdMGRa5OC87y99
L8DghdburBC3Ny1n/JXPV482gjlImaDEofEVSjdMLdwt11/0dmRpuBnyxoPgakin
/WBq7T3n4YsYtCuBZhxBIlkj6UquiJfahO9i/dGfWqedUTE3r42/x9ver54oOzcH
1hbSqQlZf+NVMqdOFzVS36QdWvOlVd5dnxVhCHN0rmJLc5zZ/IyZylZOIdfolXIL
obieZx3hNpO3ahrD7lSRFHR9I+6TPOWeQJCAw8pgN+6H5X2Sgx8H84cyUk0CTL03
EJwjc9Prk8+7hZ++Zu4QRXnvPaGCQF2Bc5rn7jjhIgF0jxoFCMN6lq3gfXKV2S/t
ctjv5oTbaPIZHF+SVLlWYPRx28pcNqvBRd5hYTOn7jY62dzza+UdLt9QNImKnqZX
ZLgEnaKyHUQfj5+Z5AllwKS4+xNu/3afsv7kQe3N+x/l7cldAnaDoc2TpYIfva7X
V4FmXoPLwzZU7esJQHEY2cLrPsdmQTAOUmJCZjY6uW1a9/aqhUAhqHavBsudqeoG
J0zNthYEAgwl7w24wsjx5TSmnYTP0Z7OQvu3uZ36LYGaHRyH61D2IFgyo8wAXyGp
FpRqCE8APNkRwqmjMziDxgNj0dFu4A6/0Wi9MxVZ3yxnQP7GrdDdsfmAxshGEmgF
I1jIA9eUoH+OF7Lit2c3gA5qoE5davaJZ9GQmPzZJtJzImCdIGyiY5y+T7eBdQ8+
KSBPPbAF2ErkidBPK/f+d8hiP1I0eu5zj2FGk+yGWVRBRSTyQrjo7Y6g0+9OtvYE
LYkQXP1pCA3P78SuDnjrgOpk013GczkD9XVVKPXfYxb6yVDQteuBDgL+6k8CZhHS
c7y01lXtFK57mRDlbrxn5hB6gH7z4WYmkFTOucUlXsKr7+3+AjF7wjLL/UQWCE7M
64uTwGTN1gaP1/hPxVE/fi0jumt9+A8OeuPFUEV1mxioniyFnaMt1j/nZ5S8JAXM
+IWFme/PgxLwfakQZDgWnxVseOBRVZys9SNhJ4YhN3HuxxKb/yLQ8w/7fF56FWQD
+uX8pVTDJXSLne1i6NFwnMKLSUIi1ylpric3E2EOnyuPAaKVJ2oFPalytH+O8a2T
2yFgaFCz0PC2WvLlG4sa7xnhDdfDCF76k/6EC3wi+yBGZxdHAqf+H9WaPXSFBQYP
rqFH6Uq6AJ6y6wIVWcsvV2zn0UC6Ig/Ie1qwyEzVJPH01RP+9MqhPxSICQVJmOz1
yAsjvdckjPSZmg3uXmNwKAn9IgIi7X4rAg25/7zsDXQu2vWRPB3t2EouX2+mRFGT
4vNBYTVbuFTqkfVluy4qaQOkj74lwRdCuX9qb8kif9H9+3Njmkvy6EDiaX7wxwT4
cOOaSVq4vOriKMPzufz9qcIEZ1rlVYOAdpnrfrb17RRu0vezb/hjIs5B8ayIAMBY
OKYaF95U+TKQ5Hl3/yZliYjPhlFeWQSvi+sGGxDfVDHThPHJBPjkmd/n7nmH8UtV
VFq1ZwaCUfFGmCp/cgmJn/Q854GU3tEkbYOF3LLygklp/7OhYSotdwKFz2HG7K86
Se5cI4Njxdwdgx2KwMNMiezNu6xvnJwuUKULlDqXzkLAFYzHy2AP3qkRicTgIjYj
DRlXsD0ouuHl8noKlBYRmJo6P8v35x3uLJezwgLIAsBJNNYC7tHktWIGDFNdUUvV
Tu606bgb7Owbx9ISILPkR4vVZJMi0b2Jmw8eg38QLdmIfqTPxnG7NOfQFcCzZI+T
UAwmlBFWY+Z4a7wCYXfBo08RzMWTN+kbjA96ysoypAPo7Y/Vzy5k2pUf2t72x98B
ngrn65ZuA+JH4/95r0ZB4CvB4YfhDgDuJfa40l9LWRJNcj96hM1jdELBxT4f/gOI
5gVGzdKn1hP/k2CE/XVJ5HB1RBY8BIJsbcy3S4ADNrqirj1ok9mG36W2AfRzyCn1
7jiT64R+qqHva5n9pMSx5xz+oCk3e5PkXH2iyYRV+eboUybBis6mSb2yEvjmDBrS
8jfV73hhREDNddzODUnQVBELx1BiEu4f83A39zpI64bp+o8izQRmBri2/5hhkSan
y9QJjjUguBkXpFuDGHuxIrkdOKpEmPtoTVu2JYlKRd0dz6+JKTH1DNRAWxPduZme
Rlk58f9HouP1ZGU/UBp/QHiopDV0u+IEyC6YbY3SLQQsEWoOdZqGdnplmhPLlEaj
SRika3qBj1+5nmrlrCgVKPEAYEDo/1O1IhOvWwX03I06HQlF/jSsrlpzIphcOI5L
4PnaLYOl6/s7YojcdS1wyvU9nVN76BNCAyx0bXY5OaRrk5t5ljHYvXtzf+gg1AHN
FtIQj3yAFWSUjy95ifhC6cj5AYTbXhXSw0gR7EtZKrJgNfooj2wS4Ahra9wmWrwA
3QAPq2uXq6l0P22FD9js4IcU/BHwACCjyVjboQDTj70jF7UKQMmff16bRWiYQxSs
+/wus4jiI71q7Evh9L9TfDyViUrucXMVBL0uFUvJ4J3cSsm3dKKkGkD9JOx+IazD
iOeND0ZRzdRE1P/VozuY5CDN4uB6m81gk/eoghrf4BnZR85/WkScbdcMli0LSDK2
H4w/7LDCSnnQFCbhZWj5Na+fwTVYB6ou+XRdL0B/CAeEAOkrwuIo2Qp/UFeMe0zG
rf0kRIgcEOZppIGbAFuOrnmPTNkmb6ijNMDUoJwBuMJyYXsanAUs/QpFoNBDX1QT
xqVoDVoxOci7rK1h2YeHSo+v816SWmFAUJ6Fg3wxx4a/cpIkAztyacMbJalVvn3f
fr22QgcJuWvtBcL/gGBUxltJZpRjyPVb5L4uKCqQnAX81t8nx2TxRxRGJY5Ez0z6
teVdiirjFPCuLp4dDPLj4AtqxBijLGortxbW78xOZY3W5YnkbLup5uXRwlQhfJGA
ZSIojmjFxQ1yrU+xwC7f+mg4aeZGfLXuBggbtTtxJRhGR+G1nOHuuvU1PI1e5Jk5
i1CvHbKfKPE/kauoppLt3hm5ScuVTPqhigsF2iyseGua+b8D3TvX0Q9Yy39jGCoG
pQbwOo+w5yxPy4oqCN1Dx/3FS49cHmAR6v2lkINBGJpt3O65qJWq56m3dMOaMWYO
77VAMI0B+51Hld+bSktCdluMsfFUDMlL5TA5rb04i3AjvPCepYpJNrqXLLsj3cQ4
f7EBUjpKsKwRQB/eixOhDdNYC3QZn3pxjxhgVVZcO0ybMkmStKfPifJGLutVf5BN
s1s5K4qd8+mIAgXwrxL270uAqr0R3MsKzIvkJaNf+lwP0o1aENJUqUQ63rD/bmGC
ATP82cogocdVEQYGuTJEW8wwiHJCqx9yHp6b2xWTgZjH/g3tSjH9pJL60z/S/iak
E1j4QNMjDLTxmzxbuGH5lPwcMPuXrhW1buvqR7NY4qghhOrFL5Ftl17pYq8+V3Oy
z5IyEJMmk4+NO47XM5MTSCCd88ruoF86v502AbWpj3i2wa7GXkZCneDBESjoOoV5
2U57N6GFv/JvCDdz+lX+Ak4q3Moj6OgOakKY9cbOh1IxSXCYBFJhpmaQ9Lfzlryy
f1i2wAb/Psxzbl8NOMfKX4GJU5lxeox6ms/xoCOgGyKD9IKyXTCMVs61kJt6Wi41
3NykMXAT4ewqjDo6a2443nWxAhgHOj1sLfAllQLsHeka+ySUSxqakhT785OfZZEh
fvNm12DLCYJtE9Dxxoq6j97rbd2ZRINrQE6RBsGk7eCKHm8BQ7SdWppgeLesYQaM
RroKKpMLs8sHaDLkSlmXIbHpEd3t98S0nFhFXpeBaUZ94glGlQJIbmEnVH57mSqY
YEwFCSp2bAYu1RnyWlCt7yZCGQSZRhIzkAVulFFN4Utzx9dP9+QhXxmm1NqBv1A1
554i8/PbBeAUBx7fvwhYQRSeWrWE17SYyycTZc1Mbbl7EyqF6T3ApEhiyWPpi6TW
EFvPDn0neYxjAW74KfCq9iFHVJ91YwFCxgZsq2vCC0OVOb1opVqeW2v+8I4yf3lQ
ck6qi3BV2U7tFOwEmCUVUAoRKEbpTPFz+puhkj0THUWx35ZIjgfnQW9M10ioIN3l
1IwvX0aNxFTEbcUXB1P4tqPhx3R34qZTTxZwL69gG84jrdqUozmzKVMhYDEc5WdI
U1Qzsn8SXwsz/cLTuBCju1O+oAmOAxvfSLINwpLsdTx7yjLFM7+HMRLzlyT52sd5
TdHmuh60BBGiYXdIC9k/AKWy3x5aaoTyNxlnFJOBXXH9epOcIOCSxcVViSdl5tyI
yQ2VRxT+goJgooCmGm8SpFd9/gI+QeHFmR49OHkwwgW+TRBZ/XMGoPEmrRHYXpe6
Ella6jxxLH006nWgg1mHNs2Q1W9HDA1OwpwT/qQfEwgGi9kl4A1dfK0zh9H5p4hA
X/dwXSvCLIcvEEt19lFrD9HyUKjBCXQgxkAi9qVaDVCPq7Y39Jrui+t5x9v5p7ZT
JOMS+PhPMWUU1FKhFHyzb/JmpSY14bEluQZLemGn105b0nJXNMorX0IxmWGmThUr
SFVcpUG9/pt7XTiT8SXV23CFivpP8b1eg7k2pMLXb1pSH0lnhGRprSv2/fOdSdY4
B5+7jKuh2HlE6cZ0df+jSSeFlbNyQncuYr0Vv1gE3PSsA2nen6BDvwiGPDDL83TO
DsWr0x2Qcv/y6+0igZkbSmC4ufLZw12JCW9VKzhQHoruO+vEDm4IzMWjM4OPeah5
Id13w/yXdkDm7ZUYco+o/CTPpS0jiJLkfB3C3MEv+wqZEewMGodecTFrXbGuEpTq
RqHc7NNttWmhyRCjX33wkta/0WOH88JqtDf/aHcIJUJXyncYpyfR249WjnEzulms
JlfZP1qlrdUS8RNf7vE2qt+7aLFe7owBjMLkTaDZibnBF+iTEo1XdYeqa5iLJ2v3
J+wFcnjOhH8c3Y2Fd/jKlB5xpDzZKhIYtIR2YjOpFSWGqDNq2ZEx8rCpB9lSh6FK
vuP9qXRy2kNqsHyshvY4rEfL00TPTdl7YXqexsGj8CU28ormT7dHuNPOi+WdKaCK
tIH1N7GtzJ1nBwO/rQmalcbCJFWL9pmga+sRvPUY40Zb+b3xvr5cwDIRS/jMvSSP
jK3bp6QqUwF2RFC7lkEsz8TE4LhySdjl8NQSH3WbDN5UNoGgD84u/44uGOq/lvsy
yImBAYIEjLzqmU1SD6y6KQ94ckvJ+HtmcKVKS+ufhqCXVVKfBNWyydM3JRZPQxOy
Qj7yGz14I9LUXempnvXbNgNMiaTar1FieQj79w6UhvPbbRHs9UQoaKXZWMwZEtAx
xTzf6tDalr74PamqcW/1Za3vw3VoZk6KFUntQT7c68YuxQS+F1LaocbL9rts8gAo
iGXOlcWLroyN+m2PIn1v7izl6+gCukKvjXqi9XbfJPqKzzD3QuuX57qLAklntqaI
rvTyoq9ufGZWhIHqgUeFLz9rWcCEvX4zrs1g+ZNcPnjYTNQIOkwSgbYoV2Z1cTy2
oqgvj7ROTaLi6HGpFkiEeS/YPlP3Eoq86g0J48yEyoanC8a8iKgfKai8HcPO7zRu
ojElaa5Muj2Mkv1ec2GAdlw74whCvYKijJlpCvGUp7XVygTcY3WZIt1HK3uKqDZK
5QhcViZqGCxM/0Doux0L+sTME2N5gSSFxNZqWSkIR+2Ajp3/pDo3AHbOCf4i+aUZ
yvDg9UtfGjHKUgm0s7fYiuym4UeJowg6vDFaAkd/x+Il1QFXWvm35HAWXxrYCq/H
L4SktrH0tfTYU+NxTNhQWVyjOGIW1nzCFAuKECksmCdbGOvmjHwYUB42ID8YsJyz
ysEAhok6NdVUJTPdwjHdiaXcthm1TO38XPezYLLnVz1g2wOGSdcTXYulPyebEHDl
ninkcD5nE8fcL4T6AOGI3UsGfUPjOR3V14SR99ZU3xPnmsBkCpbi7qRrJAWPGAMG
xvEoMjZ8tEoBJIKk6Sgc915WRXm8lJ+BeGPkjzCIATfX6ZSLKFcYneRUy1HTLA9E
3lh2+YyuHlYfBRQruDE70d65JZv1PG3AScXp5Ici72kc5HpB/Mz/60qrDUON8RNj
s9IJmZWxZ9sBoO/nq7N+6sFwkOsQJ80bid3sEv5Db7OkdZ5YsVuW5mERAWvXLfNw
Tff9tlHq8/WD37emQPsSy2r0ClbW/Tl5wXrcBygaIBqQDLNuNFHa+9FJybKBFeb0
prnPoJvHGR2jmhw9pu3mZhi7Rs5b45pKwmHq2YfpdwHpZd2wnwCwCimdJN7Qov8X
3Ig1CK4eEBKlPF4qgz4CQXKsU7CC1PdyHlBGgRTglQ+9rUC3NNjVlj6j02zerstG
yj5niLYTFz+poTr3GE8ty7ZfsL900DkjATTvXe9XxPEOLepMBspgSVvm+yi6IF1g
oPygIXPZKKT+SB6Zq8ONYja08oVD+w0AFfcSuz1xgRwU/xprl5FwUB7jgssW0n6y
uRyz3KP82pRgirnPjSVUzR/VOvUMA5/YLByuARzh4JZSNkrxMBslgOgfjLfZdpBv
ST4E5utwfBgcs/ycSmd/Cwp2NAkkNFeF0M09JPDwknS3lCoSp8jmyuMX0cjPX8mU
/xaSlc4JWz40sr30kBSMTpWGBeKWPlOZI18g/GSyWKhTwR44dYo+q8lCAaaB9tZO
ycpMFCGqAS1gqoXO0vHN9dVKSBuuLrc+a6/n8fcz9jd+g/0HQiJjhXuUAsENEGDD
sqb1lvsKZqUDxHtTlQKP81EGPbkOsGnxiISkfZgBZ6tNi4/Ie7HuLMWP/qZmBwbI
71BAWoMbUu4/4oGFGR4WFF5/oBNOhTRZDni3owXfwkDCkCoBsPvHrqswRjHO9eC1
6WG37DWkPrCsmp99+vKo94QHXJQPNNiHwrqHKF5+7MT6CAZvV48llVPZXuPX/WfB
Tk3Eu6DUBZzS1KdQoiY/feXFRGYMijnV7LnUAWRag2KdpmD2HkBjTNxz7PlF7mUn
gTWiLbJtwRNHJuY1Cnb8IpgjiTGzf76fb/RsStGyF3gcllsSd0Laj0c7G5wwijTq
UQw2+P4MR6unrWdl7PTWF9nKbNzpsuZSb2V/uPC4NMWp6g0O6sczVTgGKzY79HV9
faFnpyuxq84N7DK4CJ2SEmWH9PnoXUI6lQiXbLXf22PlWkh8wM0cf3WPp7pEg8Pc
O/sDJisb2AHK5XkABK4M7xgv5v6FnO2XKZIv2JfYYHrT9m28XCWqUNBUnlKSVeHQ
ZHznt4uLVDjoXnJgCRTpF+RnBiN5j6AOUFwSlk7qoQ8sXKIlaFPl+0LffkH/S8R2
m6c9XXTudq26YWzFirZbyRQG7hPlvh1U3qJkE2Pr0+Z/S7RIdWL7norPP/e8Uh7e
sSDVivqdJZC7dAfoFvVt8XRwaNIIZOYvfJ6v4WcpSQoHiNSpwJ9mH5UFs9s1VV2S
GREK28kfnO9efQ5JL/VuiLEaGaYI0h27ct9KjIZLuPtLCPkShf530p+RtSbGSgE+
DonvetL9r/RMXT38psPO6vtYzJ++wa3RoehjHZlSQJemerG6EsO8ZGskz0DzQkar
9eWRKG5a/6JVaUVYkNsfX627RE4RC6gUJvAXJmzP2zNUEIDKP2RUq2OQtBZSTudA
dEO5nUQ8KQzd1bVDDbgfTSsDU61nYmV2NVe3Z7USEXEabZ+SIcs2OQkWXMcviKc6
GLq0aMzs0XkoLtUIV1z/W/VLjIVyOKA74MhryBiHCdAfGsVHt1JvU5V8GrKl/FHZ
umos0z8m86Ow+xFzuSQy+i1X+opfE12aJxv8m3TCnNo+pGYGZNqmPxtCWWNlZbTI
CaYlWefPf5ywUX+mUOaN4ClitBaaWzD3XwSfeWphGe4hAy5uH+FaBpO6UUz1Pe+4
1eJFzBzUUefcsHIrTNmFD1VI7qdW5khpLdg1pH11ta6suGdOg9kl1hhSfA4EZFt1
DphRXFS4cx2B6VPajLg/AGQH/HpSCvFnL20N7ls6FMDHDTTfW6Os5XhKqJ9jGlza
hSE17phn3Mpp5NUuI261UPz1g9A7EtlsyUo1VQkeOJr3otK3+urr2iU11RVcgkYD
lFp8UGU/rURir7UtDVothgjeGwXFAwvCvEx4gIyfPEwbenxB17GZiGh2D8yQZri3
Bv0yrLzA0KPj8YudYsTjqzA5XCVsEMdOjfsbUK6Viqt7H8kIWcak4z7YbuWKDOpi
NbD15pjWDCxQal8WZYq4mEkQV4iIMd7HDXdkyLJFBTHFPX4Te48kZgyiSEyXLgw5
WKZIBbaaD64839fnK3ys+SRdmJCPXCVssgqUF3jR/qvYhLT8N/MD8QlBKGljxwYF
a/llnfL49pzDiMb0ifEmCl9JCTGYruy0yPnGuhq10+4dwI4/gLT6xVl1DcLguB/n
uMWaNIt86C71bOzzg/UgiGuq7yjxuO5itX+rlaxMkzDm/fcB9deG8zl1SwstqbnX
EUB8UEYw/nU73j/AinQYNWoyvWO4sJwnBdpC051XGi8jMIQClhuJG4OaC/Sx1K/K
HliOb6c45dHFPeR0VGyHg/P3SI4Jg/KSa7JGX9KjQ1DKmgR6QCogAXdqq0gduope
YmtBTsaRa8gxDxrPwAn/EPZ3+Jmechod18BPiX1dDYntsbjg+urwja85Ilsd+nE8
l9dmuW3yliGeMRh22N4RNjmwuj5cSYrmlQW0Z6Dmn4jw+Yx/77uv/WZg6g8CCLOZ
I1/5jc1JZaudZBn/cXS5pk9/461LUspqvr83A0yeOE1etNI1Jwh9SyyrKeDUQXIP
z1mIqJHeNiArGUsAz0LXOnzIS9cEQmA7sPw/JF1AXBak6IjnrH9qmJ4NUuSSHRfa
/izTK39lwkY9MgE7PNNbD4widlQKGI9GOLZhicrj3XdqxyY1rm1l/G9dIMAWFq+n
cuKiFYvq/u2jqeSuEQMFty2Ek/MGlNTCaTlWhLA5pBzxgWinuGcBiTmlHxiCL8Nw
6N186R59r7TZIBUiA1zIuMzXiqKHEbs+2BdctWFf+IJ8qmcQmVKS81GSOZFY2ptz
gUwAmvI+cvToBw1BAZTm4P9IBtw/GKVL8o4Iged7+cF+EHbB11voKKFcnOh9+Hlc
n5xvIAbC1Ngkl09G5Y43c/dfN57V7Nqj2SMx4UkIVk9VHoHHNVEMJHBhxZe9w/6o
RdnmUvDjS8I//jIj+rA2lF0p3TsIoU6vPJLoplis0Hjkysd5FxIvU8rHum2CM4Nt
lSkUtkR5/j3v9mrMplXXMt0UKZGCFQEbzWuZJnEdQUcbEoXOABim658VwIeJZ4ub
/wDIZeT33H9/mcD4k/Ld4aw6cNTUXCtFrogSjAbMMTlJK5yC37agSuvlQXBhk6X7
3NSdEV/bqWntUCs79OxQ7Id9XZR+hlJiDx92YsCC8h6yUj7OWtflE80LaPkEAYOn
FDU3aClNWLRseFFcw+bfNRu8qo8KebhPmTUgDUsKDKMo+vNm7iApIQrYXbbXEbrk
/68mRtPMJUfxo/nU+oPxGm/ZAlzLKwrFvbKeQHx7lMzouNhXUl0kfH2OhSc7vvCo
0QGlxmOxU7jh9quOisRoTSlTnTrFDmPkvPkO6fGekpzD2Sp7/kp0mUySsm0hfao7
cUXEDpA5g59PCp8hl0JvcliqDB9VxCMutX2feriCl8VAzvSRkoisWBlQ+nFpCeb9
82XM3Xc4JyF5puNq8HvxmldtXxOQya/g6zrw/v0ZXSb2HnYoGS+zr81pYFK4wG5X
ONnR+mCra0fYycusYoCQv0TbOMkW5Y8xP4apv9d+IToAPb/pHnCE3dYic/qGgOVz
gnTCtkUBTaE0qAEfn9p1nw1iAs2QymwqRyQUI4SvlYs3pLn/qlDbpTrxe9NcNwF8
bHuV75w21AWTSnz7j5s8oip+fBtF3ZDM1WO1BcA/+NqZE4LAOq6fv422z2yblruU
IhmfPKnAmPkuFCSSSQvgy/bTWvmSAEGPVWC2Ne6DmccREof0f54ePcQaPbEcufvS
xvIvDSBtBYUmKVPqULSVDWWvnNNiVbLpOpjw4GDBWgx8bnz+Y5g0TseLQtb/GJRN
n3byTFhv1fjaetFt7fghhdQ0XeAly0GDZjyUkmtraQdo0feoyslkxOkfGRcCSwq1
dia+wAm+xAupA1w7Mp8zMMi50OfAeCwbDFqM3C7/DEopKTQRxGK4gfNCt9Oi8qdA
odW+SP3ku/yifKQmeaW9MjGSBB/R9GirAw/pVcRbRWemeJXK1BT0ecOzGQukmueD
2EUS/ef4RTXcZMX4SMVD4BZP6pE35BSQotA0ZgZ5/+kbga6QSOQqV7gaxmLDIO8/
lI6FdgucdzE5APLW/6SOrmAwAGfSQ5BFBuZRsWONN82w+hypkAxE0ArLZ4nG5quA
MslNp0uSY1apqV+xlMMhUY4PD5D4ceZ5kSwQrIu+W7QHBeNlLEMaJ+53kxCbahO7
gjA4ljS74810Skumln2QfROVbbKTp0FlyQXfpPAjtqN25FywZTOK6UisZJWXnI42
8Hi/YkG3cvSGmbd8ARvZaoYmTw2JL09TGz/FDDaY7iPpMPOYKoWlXvWyi+I/Z2dl
rWYFbEpwYl4QIV9QeOg+Ml0wKsJ8K4/GrkTJVeyMXMSoi2St3pWv/dIcE6jIV1wx
pzx20Yg3GrdAmFDOCwYc3S3V0b9+VfGYmFX8B+zpQcR86FAeQgPaqUA1usTlQV8f
BpqfgtJb1pc69+dY1OFjPqQSkpsrcdCM6X7L5wmhMzjbGMCb3dcdc4G29k7zZyel
++nW4W6gA3+bRf6IvzAZii8llaXEIc/vZLy3N4wWIHF9/6TmSTSSqxLm/ovfBTtX
dGMUrskKBeHFixYyDzlAgl6J9Ud3iVK5ZuAgOmY5Tenj/VfyaQlMiTxwa3VzKoyM
tk/GC6vzlheQvFn5RDaQFgk6WFHn5jjQ/8eWy7xSDPM2E4vB9iLpDrD1lBqdrfFd
WvdhBdpd4ejVYV8Cm7SS9K81TU9+NGRONZQ+5KOLM3OdxbitW88xx/BoBfeAH+9B
0KNSJqNEmAmKZIPzFV6rt8x+2ky8B2QkUdvy0g8WgT9iskWcBmniOT6QKC+nWt7E
wx6CxdczedY0bcR7srML5NJ1Ei4XZG78Ie8cuI+kSfoXe0CdAuOx5ByEaVPl17WZ
v65hA3w1H4iJsNuvD79gJoZa9g1ycsWsOv6hqeaMwFvGthHSaeu9xmorgBwx/H3p
DNC6y3xh3E9fS/LcVTTz4yS8xEX21/8/9ze+G0XmYa69X2gfMdvWgELYyUhu+RpJ
jjSozYxjckEBNvHQuh6w9NXKYDWkURGh4aqJomVh43LEsTtav6MIrK2et0EueW0m
xU23iOEwBaua7QOOmQk/sstmEqQP6v1iYLACZ7WX1YbkCLwA6cCpkGMIVxbaKHf6
DTzoHWxaACbrLCZmrM1m/sIjP844UxxH9eZobuNV+p8g30Fwlg+KSSyMse4KS60L
LwqMGwWaTQiSIpClRjOdqhSifPyQwLYWx3O/TGuQN9nIZiW8WAFlxAJulir/N0rH
h8eFDAO9ktoH+Za4DFXJR4Cfzx4/Dqg8iqK0P1yumidAhwLRoV76miPk9teDaALz
VJ+tSKSZivOMEwa30OloHj22B9AbRxl3SwDvhxf2Ix0WnnJf2UwXHZ9jovnwNM+X
XQAT4Oxdrb/3XjHZWhWp20qKU09VrGxx5lAmhauoGW+V9uhlQ4Ae5+6I7wiMgJ6P
Fsr/YiuzE7tlgJxFAeVQcdq+3Sd81hrFjABDOHYpBMNZTQ/TnF9QP/KWMxFvpoek
WBHvc3onOrsiXyxRSFOvaFWXpHDuva0PkINA6eXpvlm5R+TuxrLLLgLnVonf0WWP
H3TDug93iO7TAAlf76go8wuhp/Kxz8T5/gqx2MqmXrFwOj7Ry5y32SsbfeHFpmNt
gpYezoccJi2tDVNjmr8dHXJu6FZ18zUzaN1oWGkZJLn3moAQ6v96Q6NzrDUQDRgg
bp3L6KJHZpcSL1DaB1Gk49opHHbWYlpFNM9yxDWWxJRnkYvFNfi4+3BVzQw5JXqf
FdrqdFYtAvdBjZllWLEF5eaBwm3Hl5ND5HdJ51VJWpru0eCLeGm/mXDN8FSmhwEv
ydVqtcyI9yrIIYapt6h30bgLo0kbY3YHb0W4t+KbWidLxkVwSG3/vXxwpO526XBF
5DyyfKdeuVNNMpio1jRpCSoQIiK7eNrWU4pN+oCddyh0GaPmu4cmnGV2NOLqsI84
eGCw856UxSV0Vz/tY0aKyF/t5UVJrSj11Fwz5S++cyHkC1zOXfBD/O6DmzvMwS72
dGN5Q0mT+qiFlNUWo6UCY9t9nm7fjZC5BV8edlyhODdHW/PyI2tmbe63f+W5ut10
sgUvVmxMqaMF6t6KWfS0H0/vIy0D76v/wZP2YMf9LBlGu2JyM6rj9LvtnFELD9Mi
OyC2jZwukk33o05Ec198DcGHl+EuJnRbWH6SGpp7yCOG2Ij/uqgBnsvqoJqCcDLX
3uxRefvMHTfjk6QEtpGQFYut6jhd7Gr1cbQ5jrlJeiYXXOwxzkBhDe5/eqF7nGne
k8bBw7DgchmSQ29Yi2/xfEWQ3j4gC20Skke3TgyWQ/7x6TOa+GlqBf1M0b4g4PZo
lAysbp3aLiw+QoOKBqIrTq13OSiB39f65DpxoTWcBNk3wH5uUwhaB4jw1Xc0B39L
UlVwKTbglxz/dFkdiRz/0isrGLfsaNTYaWBU6DNzN18ebRLJlMEz0Pmsc3rbIr/f
capLSNYiawUDhEOn7vc3DvXF0IoFIOA1HQWQhCSnzTHY/BYsmsBWEPN+uuK1Qom4
vNhdrw51UPBhd3oRPfhJVF9Qnlas32pRUGoQ1BjQsZuO0CeygyzoKU49SYs0SEzu
zYbYT2pRgvfbVQp6KA/0bYYZ1zOs/jDzszmAMtuFA8MY0FCx3QER53KA4expG7Jv
bg+gm/q1FiDBIcevpgA7TL4nZejKAO6qoD8bj+oAXhJumrhY4Dg41OBqc2ceI97B
/tW0wxC3a0MrnkRWy9DGuhIbIjjNAEmZc/q+f0mvAjskGx+NQyPn+gqBOl9jNHjj
2iOyJA815iwaNSUj2PHAtT2deuec86cBtyUCUG+OWcWpy/eGqnUSNHQOH5aTt3Wc
VHVdEtcd9kaIYL4ydQC6fwKtSX4cEvwaDVEVisMhmH5L3B6UrZJM4VvxPkYQD3IC
k1HxeqqVcm81umbIHR27nmiElh1UpfeDDRU/O03OYRrGdgtzkY3A2FKhWQmENgdy
uqF/M9zJObZKTT3O2DQ0u3LhEch+p3tFaiGxXeKSGuKwNPAztVqiDEEL715APXxl
esW9pzHhdydkVtpqc7o+IK4yhN6Vs8KuHCSF8iK9BgexR6KnkXkx353F+5KF74Fj
injCzKpevfRY3rzIQXkMDPtqjoChXWt1BSBpbI9ap+Llo5OZaqlTUz0OEq3Bbm1C
9N4G9r3wfHmXokUbUrCTTREGR/F9M4bM5mEtwTbCHGm+lKBUXsM0HPAD2cX5HMvo
ajQxipo00a7SDAJODXwgk4Eb6lfYPqcXsySdRQ+1EglzpVasFd3Oo0aD6EXGgsWt
w5uf7fqMl8tWyjREiq48/fQDdYiZ1JBYIR48oM9mFZjgfRE1jIOV1ULJN0DQsPTt
ydtyV/TdtISX/6C5zUw/xIeqlX1mhYQfJR6aVtXoWxsa0VPolEMI6brY0cnfvnH4
GD0ryvZNGEtIzFECPkGoaNkqIqVqrIaLYPAlZvYQpz/N0QZRL97vHUvyy0+9lupH
uXQvtwx2jQuq7nImyCpLpV7U4riUhiIVCOVFyj0imDHNntEhLO6J1N5Wwu1I3vKm
MbIJcAeKBPXWaOGzGWqOAlHr7i/QMel7Lv7sxmi2IAB8t3DervPU3goQCtSuuX/Q
n/f3/w+wd6dWiozIe6Ml6g0PGcTpn7qlr6a1gdQThsr17ePzMNxkRhY2bEXQ6Bho
SgxcMbVo8WwMr2T8XgKeTIinerFZcx5t/M7k7F0ncxZB6W+zYFfQm6t0w6XLIV3H
A3RpEAqpj5ihyH5u+Is8p+wJIgTkhC79e28IX4x3PzBJF6/Siv02ctUhsvex2hbp
TdqHDAspHRKZc2g2wp8ZvPhHJD0IZE701K42DItsOsywk1JRwOPqQIG0W/cgYV+v
iMH+eOg9AFhWuzLNinjbgMOvKf6XWLD8/eHpQ5dAK9ocY2DBSd9EvukSBZUS5R7A
HeDoLXZ+5/F2H7dGG1ihsZW69FVHV6vZJv+zLUp9mKPjuP5IaAgW0m+usnEU4WFO
RXV3t2d3S8ZsRHuHyDQAfmdGfdT/iQIvFBXqMO9bzc/bj+o6vKE6lpgCcLmzxDtb
GBxXD8eF+EbGwGYWRZiOML2ccRHZIk0sRtwxPpyf8JnHm53Ivczq2kWPBM5107Kw
dX5bIPr4B09Z5jGDckfiRr9YbVfUZgMqW4A+paUcGc+dhtWP5/c6utSmNncJMP7Q
qrpaBoizgzqMU/vT84CHQpqGWNQtT0rnNlhAzW3oJmz6vBTQx8aC5WWN+qa+2uh7
JMNtqSShZ9Qhk6XtUoXCINohgAcLpEGGSjxCkcT9Kbj+Yg5UzGSDDakPPAGp81A1
aI2Jy0bLqj5NHP5YHQ7p3om7ugyaqr1I3pin44b+HAUH4c4HxH0KIz7U3N6iOOqH
4FDdBFQX6EPfrjChxh/l+Es7VbTyTIwQNJ+LgSfq3/ZO6md02y4W2VB/KaOi9gv/
HEIZggIzYqf/To6nWQQTFPm3zBuMAt3+4hIcdulWT93R2EGekRtWMzlsIlGLT4OE
tB3gbQD6TlkcmBlj8dVNAJ9nkKM91L8bXOWs9y2TbnBVyrAd1aUA0l09CTxrgPa6
gj2kuOOhQIRnDXrScgybSSMCiDPD9kkoG3apm4F8zHDBoQVuOAu0MVeSoHFjvFcj
9Y7wOttU5kvjkxF5bDUbUGAdesSYtfBQjv93xV/7mSdVK8D6eejtVwOXz/tJr6Do
MdEJOng4vVyjOIXVjjAuiY7Imm8FGe3bo1rOuRfzAD+9L2YGallOe3WLt3iYkWbs
il/2UzDqAs19+ML6RGJFBypT1Vvm9OIlLzyvK664f6OanknjDzpngKqaTVo1Z+cv
Gv/uQ6e5rmyPZQHg7JvzRPlMSaQ0uIwRVuwyto0t/EkRkVmAuurOL7maAq4Z2L7f
i09Cgno9ig0d2wEWPssPu+8i6bNvvuOzFb7b8RYiLazhnWMGifaWwhXGIyhguuGz
PNwiwd+tKYafLjIydPiOPnqZ1qQbXvsuk9M7g9BK7LFg7Axdl+Fs1oAN6P0Bsjm3
ejM7M5HIaLXPLM+8z3V4UJZs3tJqY6Sk1P0GJHjnXwX9HY8uy02BpXQl+pBnJBwN
Kt1gFjK5IBYd1f3KUj4z38esDW7T4ktprDuo/IZJhGozMlD6KtpkTZBmO1K1Wm2h
TPbES6rXP1x3HCkKdzz88ljOUfeY4YvsgWuAAcZmmWu+P/pH0zRRrKR+rov5r83Z
Iut3Oju0oHYalm7DwpUAOwHmHJdSZpFHQFbQ9oYfo+WLG2txlxWC685jPFZwEOYg
aDNfsBR0vRJx5JsaxTykEhfqQ7DFSMKcskIwlkp5zHQnw9ZyHHOGsFpHHDGYxw97
ryTI8YIYUL8HfBq2EEc0Yero2O2LdkYKSZDZNOLChrcs8EFI5v5IhUvOmoVmHv73
RtAuyzRQ1b4MGq5wNPY0nNUdTOAF9+e1PbO+n72zPJhjuDjZZ9D/uHPExa87NxgD
fdYohoLY5zVKpxwuGxCOZzqUBksiTExbF897X5glO7vJVFShA2ph12fVcKkErpTA
PS/k/Jl0XU1Ls/8XDYMqngCKecL6oSH6v7QKbOl2Ea+xO3ZQ/SJCup+ISLd64F/f
IspZlnQzhMNihOuZi2T0YNFazH2ACQOdoHkO/ASwbZknjtgYPTFlYkaoQF1P3hm2
zUuaKNP3oYae4jZdZSGcqIfoMU15XQmbusxRdROiadeWTrpXndQC6g11aT1cRL/X
zPNoK08UWPc3KXDUe8SRHE2gJlaxgBWpjKlzTImEF30+6kdfX6Ot8RIyST4L0pMm
LZ4RM9sr6pt3gKVIK8ZkZTzhOaiPU6B9AZW6usgVGosfpR4fgA/w+YLTV6mh9yl9
DJsKBwUHHVIjeqiYZwjsW7ClWBX2yrr/DUKLcRVYY0/1rsTa5uoUhiFR9RZzja0J
5MxdNLs2aD7GSMvcblp/TLppPPJSLEwLhLTvdlYe4cxEM+cluohURVvMbjt6+RCs
NBwMY+n1mEj93RVoqUxt5arpVCs+M7841DhQPu+Pjs6ndAilxZUUhoufp4BD4DHC
UT9NCbtk7LC28aOQOTiAxJ+y/kixT5yqmmzGFZAHw4EkQGpYzguFMYwwYzucVary
f8cHE9RkbGjlK12Afoyza2rAkv5fdlIWTVqG93szkt2qnQcKQPY6CEKqpv/HgZbs
A3Z7rPRz0N7Jbeb3fkfND3/4y+jBQ9MKAhB/UriFVeJ3TXf5vlSbNBOOZx2NKKJr
9+TXgabHZcGc3WaaB0tIcmB0dI7mcMhJ6T87vd17bZDsEjlp2xI3J9EDBOFiks6/
SVm3VTDrWDNGjiuyIXQu7OhUB4GX1tVkL6P9rdpxmiEd0gZs1sLkwSUdgbqRcEeG
A91xrSpPUTAEIMKz701z/aRO/SaIag66GISt782WPIvrqqWfUk3sEjHHSNLqBnyG
cDuqb924wrRSG+NPz7fsamKdilvJHCN0QjlC24Upi8/+oDQMFdqoMdDYPR1OPPHO
0fn4WDrA54tq5e7etFDKoil8/C2Nnm3LE9FJyukeF2Sng5ie+uVCAl4cA7RTeHIs
YInrHE3Ty4oL4qNjscF8md9bZF93EGrY28y8WvJ6c3d4b50R53KUcHVdGR2DwBZB
6O0Lu9c8ZzAU2tW7EwQBOftQRvotev1rql/oV2muh4XsEDXpV7VlZxvhN1PB3Bp5
RcdYltyPDwLV1wEogJ3Tdi+Ka0r1SoyQgzlC42ZFqBh+Ve6jCDexXicpFdSJsuG+
S2fdP4Ev2zySdx2VzL+cQx5de42pBTkGCKqh6x/exK4ETCmDrDQZB8K7fbT2bfn4
0Zfen8SL0aHCbD+ZPhUG0ax7H31TPCRvheLfOdQfXDGbUCKFBMuPS51J9e8eeQ29
YkefWrP+QNHQfaNjAjNf9dgm0jV+MEAoWDued3X/a9iKyWNcJ4Xzizn6xl/5cC78
K0XM/ljs8+JwxunOyBZnKkWraoVi/T8qoqmkr1ezIPbwobfs+RZVjpypd/ZEPwef
oy9L8PLlTbhsoH6/2oeRijzTLyd/9A6R3VCcLW/6Uv1FDTgUXa/VTloGiIzOjYuy
8k3t3ug+WpXsp/EzNWRf78gPXjmOAyogDMJUtREbL13MJpd4y/U40QRV4698Add+
/b8tkZPJ9HmL/lF5YD4N0Av2ds4VPuUWH+Bk22ZlXttqdH1LBmuULJj5KktS7rnp
YgC+QGLvqpjqDVX+f8tG27ob44DkkGCy0CxIAC5t3G4jf+dWOGUd6b+HNdnolWOn
IeSZDf9Y+TWCSuSIwqNZpNDiTP+wjpBh8KVvGLle296D3kxnECRe54UgiI9CBkn3
Y9nUTuaCF+HTcpTUHirdG98nsMoLy/1pxcbfrnroMeF6iNEpW7N/aG7fyeMdOZKz
uwhw0jyabs7COEQSExfksBsIP7uhXkYuWD+4vFGbk4Z9acRmTjKnW5DIHkmiKsMW
wi21DpIYOjMWdEXrQVYwNcauNiVrsDz+teQY3yXXYRBCD9fGb2fYBjfKgThxLxvq
bxFZU/d0rKd7zB+utnJItYvgyeGZg6MRiy+CN4tAsjOE99dpMU9HpBPDzQP4Zy15
StLQ2W48uhSjJIfEeQapy/Zx4UZRS54hr3n5h+wOpDZdD2D7vDsx9KaAzxHJ55Ct
YRhyYfDx5qpL15fh2eY1T1B7l3AG0uX+t0YkvetvqkF0Y90IdSNw/cFpGEszZpSi
GwR+ocUxjI7WoIDZ6Dq4aTmXBF/siuCK/chHeaTwPaZQmgpOCYL63Irfimyc9oMR
s6/AfUeBkcuR1IFq78c5uoVVFr6TB3abH58AQr+1YGZXc6fJuCj2Ea7e2yvxKIzN
QjQ05wQgzIF3PuxufegZjHt6hUKrru3P3endLvkwhaTdOPe1RxqsyFkBpzoew+ZI
ZfuA0y1c/jh19eBOi4LsqQW93j7nrH0xsXeFIAup9Rr0fJxUQsEbH7M57cvrZuiK
i0eHITz1BkKV36jgTH8gHW50DMcF/idDplwgisVOGBcD8iFRuUhXdU6W6+oU9XP1
tHdhQnaoIaZ9W3Wsjpoh/EninHwDlh4n8BJoaFXlHyTkZESjXGcEd3kxJQtHqASg
z6vV0XGTmi3aGlggHyJwSeRZNs8h9MfWi5Y0dNrG5BTh5NoD8r38f3rsBY0yIf6Q
tQEVRBrHCSXxfWIQ2Y854KwXjMFIeWdJL21cFyt1JbR/ZwNdrhStBgLjAHCjIQA/
lmtYFBPh//6LyvhqK+kWiImZmJT1hKY7uovw6/MHds7cZHeXZwV/ogBbpYwX1vKw
q08DCxB1u0b4XY8fC+AMzRvG669dD7X3W/4nxEeml+orua89fufgwTPwrrPzXETM
w+/MG9dgqSGh9WsXydoENkca9MSBHNA8DGeXiszGSyql2h/06bA5ax7VEr/L7KU6
/hzK9G9ACB5oOo/k8CqRTIIcWB+2ewzdAlwrAozCyr6tLTUoYZimmT+5F+Zxn/iK
KMNRYt5ki+ynkn41scbVQETRCwL473ZxG09Si4d5izAblUnP2gj8hu+0Y9Dtd0FJ
BuVB7vMWvRlhPmMLM8Fm/iimKAquQbS3htnI3cCAtOJoU3xCGiL30thA/Pk7sefQ
6pUimMTku6P8PR60ehF8SwxtRdUZcKyOT+cGm4P6n/tuMbfD1QitfB1ypvRqNRhy
iKS+VKNwF/vjeMKXEl7sWlYdeMjUeXP1aTb8jbNiz7GDkHiGqDjAfsrAhI2n7nty
PUa+DDfocLpM5PZa/Qo/uh3G8/QaYdbxMHsvDQYfxvN8lBDv+4Oyu2ISO5D8X1fV
xO/TqmiJEjMCwN+ZRWjuZtEvfYaU1CR+eua/rBMrUVFpCKJi+0TIg4zehOUraOCD
v59Fe66ILZxZGVg9TXlUn1jrgAMxXtSJ5plSyoV2VQLDYlOqDOzPtlEq40veFaIE
FjpP4q3vhAqeZuejRYWqJsCZ1GJN6OIuxUWV9ob/zbtRsZcB6ZQvPEJm6DM3JrYS
nv06F28uVI+TC22AXQ4c9sd881VbH/u8JRxnss+1bFzAnIgt3TXhkCUF3gmwBb9o
ELlBj29q7msAcZPDnqjTqUVLG23d1jC2SiMHPMoUrbiNu+QuYwugeMxi6Ee0N+/q
noi3Ah43e34KdDlfRlEEr3Efj26vzaORpaAztoDenoaIeI8sNPDu6rsW3xRp4bma
wF518lB5C9lILggST2WWkxep6qCiKhvSzogtqlKQCEfgCXm/pKrKzyrBnRjslNUY
u6Zgar79z9ytnda/FpmlWori1LleG6/vIsxljwivlD7liXJwlu4pot0ONi171iy8
82uuGAgN4ngngMtBdijTh0Zrc5s2b3YJa6mSiWiLVRFa+OQBVm+gd/QVxl4oMG2S
0WgY2r6vJQLnssRygim+Cm84EnuKnfVsKaGWxPLCaFTfAXj6fWvwKwGQ9zloXvsI
xyJu8tmeNGsTLvRwOsNvnm3umTKwX52+YKRQz6oPQxppMNkaNuWWcUAXGxxtpmVU
2dds5ukf7HiAd+m2sGKcp4ZB5fz9QJMXKaBaF0DkX/8sSzO5dn2D9UszDauVRObC
PUzebPpkmEmF7oikKUgpSZlG27KkYyvUIc/DEzNtwHmeP+c/JKDUrIXikZmSHxRY
ou69GJjJcyBFZ/BiC0+RLJO35EgdjrG6w8ASwykZ1rzLHjR1hb3Fd1tlndczAECs
4tvRvYLuMs9/h9A4rEMhdSkFWvB8qZg1eizXRw/zQyvChBR22UVzybtJLkDOZob+
zQOLL6WSfo9mxwVw7XMP6xejtTp5bgA0gMPQp3ZiJncdlHSmkDijexkBoc3U/uZX
cM6qH8J/+YRWlFLaAhSKSs6+EvmZrjUI7c1h8F1gdL3SpCq0ZBcoMJ6el5OGLjVX
Hsfrd43flvJiY8kTBoqiD8dNr8vJREmhmUIcHR0gZ7JWcsHpPa6BPR/YNwPAipv5
kDSaxie/Ii9ldPUTTqFLysKJ3H+nIzSYKBpTUH+nDEGmsP7A3PqOnWxnXjBDITj3
3rW+wT02kQhNfOCqxkz6qV1hRvpwEr8ka3AUbog3af6ez7bnbaTRoyogB0/WnOk0
3vxFZPugQY4jvYCvzvAjqrgSTeqrLMHEwJ7NxoXeVGkGgnRgLsUmj9i43U3ExcRZ
wxzI5erwQHEF8r3EGmII4WAsw7kRQAnroD6ygZcd8rjhZW13fVJNRz7r1q84COJo
R8IdcjuZWWlwsWYGJtVEaF+/XknIEOiJkFPDzBO8okkmVZ1+hDlBYJfCMgg6VYFI
4qC6IcNDtudkbnaPjOXoRvGDLGDYFN6w+91lNZA0yw84IEhdZ0TtlZklGZ234x2i
rZrqnlX8v3JBdW3UnpFxkZCLkadii1HV6WNzjxGnFhlDafmCE2DRJ+TshKLoR0L4
nBmPWUxjDHEnN7Z69x52wNQZyNqmeItbuigRjSdscjtAvPjYotwCLdchUnQxof6c
C286XefgilQjoeMRviHflGtiGaNqkTZAL1xdM8D1vBRswdeDpnUz56Q/7+yPKxqd
edaygKjU7sfAoUDADjtb5AwEjST5e5EmDo7wsKX5tNwP4LhNpHRLhy5SkX8O+ApR
ETqjuHHhhyYG3QIpiAdXfdGTiVUGQFNXQ3D4F1K1SlOzws/aDtVikv1JUbIJd01h
hkiAB4WdrRKH2OJZY4aioF0qd87IPQtFS4lXituEuv9/rxc/4/g/0t7BiA3bc8QH
1SShEJ8UKDi4FUqSMP6fpRzXgdQWLjLZOYmn3Lht2XGz0XQcVmtNTeG66xlrDyK/
n7PXIyzXEz6VSDvvEWVh8rUmbleCtcaqTUa8Ujzmdxp3qlc0PxDJmHp2cQYebBrg
5+lOTF4K+WzE8fdLLTlXclNnB2p8yRgE5QSeyPNE+hAnvtmBDRRgOwTNikXb1IHT
exiyj20h+0fP1FNkuntdOPub1PzRd4uMJQtOwZivAKDorGrtJvkz3CvWGej9BHkU
bumtM84RvVflNdLlyZajXW2sP5yQoecwKwVn5hnrVH6H0VnTfY3qICxxONMoq+PG
6ccw0WYJ8Gr/4YmyslNzsroWRm5DgVOQjM1muJ5dqrjSkcWTWtcB1z5g/c658fvr
F09A408xV1ZMHrxL03lO7BD6d4P3DhzdP8GJm37pCWUm7pi45jHZvNksi2X0ke0t
Ac0IwVnF3O026U+1eyIqKtgV1nLBs9NStfdOm38P9Sm7ZWGNJ+jzCPThQwexuxpo
mpwNyS6QmWDwsPiztAKJ58giAy3hNYNYZH6lt20/3/NWDrfXeAyOG3aEO9pgfDrq
qyC7Q9mVIsffCWkGSxe5rkrjBSvxUoBl3bdL8SSmDZ+6sjn+RKWzR/xVs9BjvOq/
XRIKnc03EYG0ClAQE+aBvg95rRJjejwvZ4v4uqVbE3D5IEkNuCbMP0BKGALJW0Ai
dzvRC+X1/imeo/jUQk83Psa7zHged9KccxabOix0tmP6KIb5ffOsYtUt7zFLIsqq
n8lek++BL964S+pz6zRNx/Fi1kZBBK5JLzafqoC+9n5IOMPXM3vrt7DudDodFpju
fyn5AuBzS1Y9lHVjZWHp9Ih5wttBy0/V2DTKeemic+ivf4PWeGi9kQ+Uh41RTXpP
OqdE+9tBsR4V9pUPEaD+Ge0rsA/gw1Iwrp2xKlCp5aPvD/yfR7tXWr8+E9BV5ivT
sV/VCv74vhTYv3dGIzi/LU5HHSxWj+xDFCDSQLa8P1/Xyv9dl1UBeW31gJXAklU6
W7jrzhaWZtQjcBNg+c/uSK8+/7ZypZei+o7AHAVWJhBdUkk8AF8DznABsIDNWVPX
58uzVSZoU/lvzaS1mxOhOxc8EVKl4MWSEm+2PsmNqx2aMchMq1Nnrbu3n+REzg9J
WWXf8D3No7F5lesKAGpi6DOrbr2WjRHA4XFSlgMoldHDLXNp/6OpZoFOqBNMdT9X
tlfidjUWGG8wLqQ2SmS6N9jjgCy2l4Jj1iBc6SIpmcgkDjowQSv0CYDDO921rO4t
mTzRNtl/7V08QT68/iCRenuz2vx+30fZGdpCW3F8mSFb7KRODxOQSRTTgD0MG0h5
LiRdjXkHYNHnywM1kfi01nFdgaPsAT63t2wsjxSI0ZmP6NYO8OpeLiHnxHPGyrVk
GbpHS1N8916mZFZFED56zfT2WROwkzE9ljnhm+NnCCn5EAgJohQwnr1GbsLIHr5i
yQ+B3NKJ6IgKSG/JlTxYcofU9eGvRoIRAYbWiPS+xS1n1XZWL1NZHT2ed5CQmg33
OcnPUIbBZPq77/kVeKf5ex1MW03STFvLJrHEWEBu5dC9MrleDl+5ulMzd5isEDb7
FtdP0fHLVe2X1noF5JS+iV91LL4ZUrtPBuIGKjgsx+beuIU0XVq2hnfKZLGcZr53
RT4/SmGq0RRqJRt+sLIPIjorNAfVvgF7TyPBKUgN5JM6kUOaqHLR4AQsOj1jIIJB
u03YGtl2lVoUjhsDux2Iy3Gc7wzjuPtaknYawzpON91H1TTuhvYUFIdih2SIq2Ae
oEZ2Ys1Ppu9VeGAC0LBop8EkLyWJQErRYextKmTpg1CkSV3QgvatHh7c1d+q4GcA
A1LUKIwQQIdvqiXxKHr7JZBpEezsHN5CsCRMp4brxN7iufUhRpxgAmGpQC5nRiy3
rzaF4e0RxBOv/DOEW96E11WEHtcE3SPh6KdPi+Q1LGTolYgfTYpjqYUnr8S3pmID
lKVfyQJPDU+XZT3Zd8Edd8U4n8CCOpKCNZatrS3493UXS5rQpCi+K5xrU4eERkA5
DLUZJNdirNCkB5z+jpdd9B0C+r9ALYpYifyUZOJG1A8KcOxBoJDM8U4cRak7rhUn
4kLPZRV8PMC0VSU4I8tHTFcUpdoV7vS/x/4bLbY6/meyOHMRoZPv4m9FtoONcAi1
Wj0uNTBatccYdsFo4HfZQvFeCg+2CestFj5TueZK1qByP/SEuuRuNCGSCKsiIMjg
LUsJUPKtE/Lh105O2iytcbIMccXCO6l0T7VGBrEULbE5PA12TH8ssn/obSgY1di0
QydcgbTlLK82xleLWKBY570/txyPZrCSSjZGrCVAb/2LnkK/BvRRkvY+/5nSdgVK
M/2dIHd7QZOfIgVqqV28NlQHVPmSqWUtpB/2k1rXjufufOzLQJ0JAi7l2cWNexYB
OU42TEtL2Mtl6M6nBD6BHRgRTzUMWcKp3GhtvaJw0dw4hYhNTvsSDhgXBFCmUGT0
Fcw17kEDfUV830r9QK32mvbK8oI9ySGxMIV2oDPqiJ7Y2ZyrzzM6nC0VUBQjdekv
BVzDXoz36biYsf8aynPwRwz2E5MA6HKhGDJxW4byWbC+h+UdFgsKzg6EbJ2CRP7U
NZEF5e9zg2FA2ubfHOXx5vAyGUJsTHPVA9qLROaPFdGR8RrIe3u15BJ9slpR7nmV
936f8MUkoM34yuN2ER/yITL8e7or6XbdVgUDTegNEZBWwBjRHO6ec6wRV3Y6V3tu
OdxaAUK2t3a+8YfKvlg7rWZWrI2j8yAw+/LnstWrV9DF2mK/5mY6c0Jqzv5HinE3
cGivvjRD25eU2czysjALUCKxm+0mfHhd5lPuiuJTTE+D2bJ4raAkqATqSmuCY9FH
PafXJ4v5PlC5o1ye/WisZkmdpIipn/4eI78Ka7ACZPTKGbMYL/z3q5IO29vL+kA7
SjX3r76F7pIZ0wTWTrkB5fgkkciRKtaVHg6YuS4eDQRDZbUgLkv+e/jfq4p6gJqK
fbIOC6PMwQIQRzn8ZU8Fd/HfkX24z3AbDc8NsCx/Zo07/uE2ozPP4la113t7hHJx
kpbMyefn93PBmowFsfxXSWeROGkLF+ERXGwi50M1+HruusHECkiCWodHeoh2UySb
wP5bh1H6Rv/gHRQIGivYISaPCy1vSkKNpcuES5pP475QRgaR6zMETMc4eYpJSkfK
HAeS8uT87RvzrvKSK183YzsTY1kRP6JHAdQSWv6U/6iVcxH19J0ukE6MQwZZU+41
1ZzwWB/Lv+JbkySbcrk/ybJRVKUJzTGeQEiYheVtoxRr7ZbO7TAcvkOpz+j78QAo
G+R7CrA5MZGVHoRp/t81xRvs9kZvqODEPXyA1zklePJvyBvv0EyopjECJzzImAR9
zKOmS00k7c5iZBNXDLndqjNQAx3YIqYR/m5/vu2S+NW0rqFEoJRgHWlyBa/w+ofq
617Er/RsDRxL+xZOv96Ip0Ysp3/i3oatuGoYSm1LJs4bE16Eh0yHCL1GeIf1i7TY
QebZLYHagdTWS5xRf4HWEg/qjOxv1xHz5cmzOl+f+wlUy3qN2WyWZGCCQWBoIuPV
FmRqJRN8+pnDBpgv3M1Q1hV1TS31WbfbUBi3K9568LDZYsbzC1zYTwq4hlcmaQq/
sEDx6AkJ76uwyBI6ystGK/dtxga/5QMhzQQ27NnEC+vXPuKXXmcXQjl09Yk9yx49
wXgKMLgGDQs0rkFDSpqfJmJ00g+EtyjjupBMVXYK/T36BAXg6fxq0Z4mpmapjtNm
9XAu/YEsbU8cCrrwuYy7e1NRSjpwzvJ6TiFkl6S68O1D5wko0pv4jwHZ/37GgnXi
k6tQ++BBRi/jbgPsrNDBnunJzASjiEPdCQWEu5IlZyIGKwKK4+i6po82nx2hIy2l
uXOv1LFFyJFGFVAWScgorUAVOEFrCy5hdndQdjwV24qLdzW9crN0+MycyWEQJLYB
96K95VevBz9MhERkXD6ZhLgtA2X9M5Tg7uQk+qY6zgRhyr6bnIs6bbnx7FkhIFwq
ionvO+yQMDsw64jNkWIWhuvLlXgTFjd34Kx4V++RgoOOBxrJDmQr6CpZULriyTGG
clhZLFqBMJ877ma3EHYG8uzMIYY6HUQ6x99fm5bNKu0R3AW5CabJ1eHEuZ0xFRN1
1K5kaqS6AykSaENv/Tt53+GR++fBG5i6FhJsjQe11v19U2EVmPRr+7Gv4YVUUONL
oLVhADQzP5FViZZLfdv9xaRWF2O7cTtZhFawaS9zp4UrWrNPAeIilEqZgaPIsCFN
zdcWVL75bmMLzf4ukdtB2E25DCnHYexn5WORTApa+sbZYpZcevr5x+wmGJaWVI9w
EfhcwIq7l37E/dJ3XK+2OYfGMNYBQYo0tXYqmQcQ92XJHL1By4RISnTH+HK7xnKn
7ZIk5u22FVEtKpu3hg3m8sFiP82b7mN/FabWuKp5pZChQ9NY/iSfGwUK5rtE+AK1
K74LQsceEsIcBoc4s0UFJnPgE/shCS7RsWPMKuHfiysJ7a8Uts2dKN7qyI9gKTJI
Im+4Z3SJPmxWAVM3DPlRXDzfjLLAusaIAzS6pBX7wQOY0AYHOaicFbpfmTXyX42X
ULPq+3vMxjRIwgD0KTC1ZxC9l1J2cG6j1w/8eXMgNWsmuc7K4+eVlFu/IM9bg88O
2fG5OhpMONCP7yUNmZsRR4g+O4KFMwgv1g+x1LU9u22IDHhDWVvhHZ/3mBHEdzFE
S9VA14D50wQL94cErjOn6+7ksbTMq5tWElLL3vTPLp/XoFFwoiCHE06xxAT6L3Pn
rT430LhBdITWZem/gwUsD42wZKu3kzT0IkO+Bv0dn1cTcqRd3UEaXW7YsW0s8Cx7
DwbYtxriJTppf0trg7sNXoKoTcI8bCLhSzW7Gfbk7dSUhB0wlYSL6+bzgh/TbKpF
j+b9hHNZwqontCsxGwTgfYzK0yoJhPklJmtcKpO5TcvyWMc3SfJfke6qxNRt5xbt
EaMgXtC1TKdryRITKUwwykQBQAiC3kBFZ3rVhrPFABRV/+LiyNhhyfalItmtxdq1
POEFO42SMCuMNQl+PPtmUTx+tEg08EDEp/bw8+cbDpVRHnd0Dx3ipnPqk6J+MB8/
BdI6bRMivqz+2+4TeP08PyQdaX4hJRAjiLqWaN9Os32c7m43wD3iQUWbktVdrNUF
7Ke23x8FHfizll/bjP69YFSHRPYBU1+iGwgpXFyogE7Hn4J/3bV2SoQmnzfZApOY
62qPSg8e2+gjI8h2+cW0jbAADn+gqn0Bw63grTMinNeuKuYBPbL/JeKk7YpuK85M
UZJ8bE0bl3CEW+OMt1WWSiY744UMZq7Yx3+1U0nCxfrr1VFjp71NjW43aUv15BMa
q6uyTyVV1bn96yaBmIh9KV0to5s6nwgKZIifsJpcOrBrAB/RAmoB/89y3RQBwq9p
CYCVtC3p/KAF8L6gXBu6mfnrz5Ed/vNGPBIkm6qflNRJx95RCnZVkEJtuJFJUe+f
t3T7l4PtxKUxSyzgwUmdr85oq09NnC416bdbVC6LAEmX1v8RH2U/9Whq2H3A1hy2
OMWW07DS4XSKc0BsIjFRotqy4+hZhSAtjCvdpu7d9uwV5ohjafKCnRSdFYeL1tJw
mPxhu3rq0ejNCB7xYzhWz2yQ4J8KJvApTUSaAPfCIWbb3tLGrMi7zol4U9Ig023Z
UB5J+Mir10sfGU9DuP/W/5Fa1+AR5p9+JCC+mkM9NA5VB+KFWRwEgRwzIwQs08Xk
kNvN61b+e3ytfUrP45Z2JSSLHrSWzDnv5mZAMAiAmGHU1XEn4RHScrVMYTftDb6p
DYmL4E1zddXf/TKInb0YwSCrIEYjST3AczLmdDgSX+QRXc6CwFiUjHo4NI2sPvTo
tM75FtX/EK1+NI3VAvhrcaqg+SLqevrPa1RwyfUDGaFs3fT1dkEGNcjSTNTqZra4
S6opFPPloImBdK21v8WN9wuah1BVKEb0DlI0J+X+PJVUtPjOkA546LyZR+zpehK4
Whhe9ebD+/s1Ys9Zj/RobTZt4JfUuGbvHOrrpAfYT6kkpNMSLfiNWgPJj+DuXDO3
A88Znf4NPogklVthSx052mEXJtUOJyFVwr4ypzCsyTepQve7FgPrI1iu4qiI7fCF
SKyJlU4U16extGdAe2dKFn9PjwmSQ5Psc/jHdWbdVUu4fxAhRT1C6HUzq5cWkvQu
1qY1eY06Y13WQBUOXxDz8QFtHg31InABm6fZtQoUHn26OVYk4yFaM9oID3dqUuCB
vUy371aquK3UDLDmo41ovWFuBDQHY1l6IIkenKWFa0vp4wYtVhRN9dVM/ue0sTaA
XMFGkFA4qm9DOpF7XiMgyqrkOpO59gheiFDa9TPdwbKMurxI76XOFgDJIrYliB3s
3IOej7DHLW1jn7kyIeeE7DywJ8W907AYCEvJIqqIETySd0QIXSa9704U+7VWX3MF
ZuYxGGSdE8M9F5Ums0CbWuUb1GwB2nbPrTyYrhdHXRL6VDPf5NN1VIJKcL2Y7X8e
sLTn6eTqA8sxMuZH3E2TWPagnbqCNJ0VdQAEpvu0RiC1c/aMfQQXtRWkWuWX6hvR
hb+hMn6/vMIeL+P/vRSp9LTo74FH4JZRKM3aJO08wbsOJBLTNtTQqH4OpPSC8hX8
WCDavLlxSdiHpWHkUfRsApFJueRykHQRdxo6UoidiO/AYAv5CF9Nm7F01SE91XIT
MP7jXggWa684ebHzNRRQ64OLjz+1Ttwnw9QBijotKY3VdUGabM6KVqVtwWOFu8Fj
Hmy+4bIvGNW/TH4xx3Pp9/mUyZ8vZENutTG/3XlStLwwFiAM4gtSbKCg+b9r0+Kc
jXEP6rFW5fjrwzQOY+f/PAIqKl3gDnVcCD0byKVN77+znDRYURp2C+Fxop3Nctqx
fsoe/mLRb+w5q8o4qov32SLt9e+UCr5W5jtPDMGItL6cn/ugfHgfi3kFm2NRz2cK
P7rrMMsBjHI+gwf6Bbbdsfr11fmNRKHIlnh733RhuYlcS2zItUVQDCHzhpwni+31
0keqOyF4+YbKpCeBCL/dhSGb/FqI1OeOYtv3PlG6+nkZveeL/6PhbdWaMQEml2ST
hg3wdHCm/gLa37Q7ZRbr9ReHQoHqQ3asgFegMUdsucKj4jVbqh99Bg8dgy+PUJjp
yeRUJRozfq7QUc5wx1atrx6T6kSPinobH54j/PFkINo25YdzKeZ9VDJ7xYgHUxcM
Hl72r/+iO046Y4FEhGBEhW+dIvuugGJLS1U5Oc0HlF3CqfRg2nPnk09MUQmIIzq0
Aup6tMzEOlZpRdRg5yKMTl8d4zt0vLwkANsGWoogDxmaaO+3IoZX/hASiKJubZrF
KF5JLXYDlAcUhlree1s7mVvSnmPzZ8oFVZ5frRCv4QZfesLLpqpTiytEQiio9F1M
lQdIWzyqIbWWMGg2c4lzgsfHGMHgL4jrOH0P62fXtZJQlLfd/7QkvUYzDHTDE1zb
P0bYHjD+XtyEKY2shqeqqOIojl6jAmfGbOKIJaTxR2QQsjYIrT19G2D3ksO0cyMZ
t2JnrmTRN6nBRh2nOl7fJaQ/YqwtQ2NC7eMS39osntiplqyY22Z8bzQydwbfC40o
ukRvHwRBY7K9OYpCC8MYuo8kneIoC2Y898b0RB3ZqHJyrmZjxgLglM9RoL8ww8cv
zXcn6YCEBmB/RG+7LIT9mEGTjJnE4YT7t5/Ai1iRdbZjBcnp5o9AABQGtC1ZMJO1
A+rOvBPpfv6vTRPApmgmaNwOg8r3SfNdrDHSTkpoRgjYSwHagcTehsK3BN9um04n
zLqIXWQkWRuRzua9u+9Sk6GaXmlCvUiVuDLMGB65T9t+axppDneOz9abqpo/KYFw
Pu1M5sBIKVkwIDC+SGhkxy+1MrAojAsbtG6FL1tIW0O70LxpYjhV5Ik63/IQ+I19
XHTwm1j9G5kMaY/WTZayCVPCNnkQvjG20AKNbqAjYGIikBpEkUqOJ20DR4RHZya9
IzSkb/tvT1m8cmE7NBJ7ocRTjBb2QD0VKm17rv08Gmlq92WGJa9Wr/gEwHCc8t2M
N9dGUKnkpNAiXNM5LAEYM0CIc6zW2A+bc2zQY3hvWE7qElcbHgQJi6sQLXnXA2ta
3UD8GOOMPl8t7Y5jB+5D+CV4zgsd17fwDES6vK0TqY1K4g6jlFhFBIuVF3fE3NFt
s0gB06ONqW6O9aiFY9y64EZEWaEYV5FVUittKeKjT7pFTQzWDh6h/XuhBIOisePA
a0jaS2GyKi1hHvtAdjZOAS+u1iUPoGHOsHldtAQzQkn5Fm/quX5SxURoqlpW7dcK
+72PZ9JxGggREfFD9IbcTF97XFEpMivReVadWJy+U2zQ9NGlvwrhhGZ0Iq+zg5Tx
OYi6GD7ucJk7D4LSa7gUUYMDLzeagp+xzT1heKD5fvIE5cRDrgAVotQJfqavg9dJ
am0Odr3GG/XiSJ62kg1r726NKoE/2bIjGQYfbeBgB5FFRsfRWm1IQ4qL0zg7LjDe
PNFv6tiRVZWqbHLnj2rq43VxhL937k/bDQ9HiSxiULveRYFOUputorT8kh5X6pLG
ulTgfcmcvtFNu7f7OqnclX9gOs+7Df73ntvuwi9lhwEenfhodwt7iXl8Dbuf4u1s
h2zoLfNtatJByzermxw9eGw8BY0CzKUytSdF8t2oR97oUK8YaLV/q863d/I41XB3
vnPXwHK7fa4K7m4JzMTEr+f9lNIGy8NQ+Xwimz8PDKuP9XCIfvSlnd6uR3LELUJY
amepnkI9zeoDNly0TPp3fANnzBBRw7e2/5HRGNjt5NvMtFIWvLeImB5r1WZKu68X
h6Z7u+JsAlCAUIWGP5h9BI0ODWH1REYIJHFJ3SDt9+QmcRiilNiPfFc19bBHf9n/
TiyqUB+hVx5vP5bFNAiiXP+jlA+3IxfJT/mzd+ejpmzDx2AxAZfvOIR9pT/llevf
GtzDZdBPjDld7xDnvCrKN7uaPddLO+x4tCFXIuarW3Vz/ZGJTqy4glAoNljCqlzX
hHpSKNRSAxY5z/9WQrSdId3BADp++yMfKxLY0UoAdD/urrbRtcvl4Sgz/UBTQewI
SPoyJFOD56dMQ0Rd4jRk5SMI6/uHP07pPju/nwG9gWiIv7S7IphV7j+ejD3jISV4
63jtl91erRgyywAtFqkmc94ObULkYKLct0NqZmPK/JPh3x7h5YjY7InMy0Wt3GQ+
vTpbTvOXvt3uBwU1fHTZgbMDIC+trkwjnr1m73+mFKZy9cajWNlhXXV6nUTrr8WW
icYwuicsa4aluJy06+jOJXyZFdUw1/Spv47N2rMW8zzeE9X4F42i8JUiNfIv0DEB
gsneEEh0do6hQTkBube/EILkQC05F6uG0mHcQGi1RWnqF/mJRfuBQq1MBvftUyEF
dXYEXbnCIlSjz2Ot8r44OGZMX9ZY3ID2UG0PjxtfLL2hYQ0tSqPYYhrRkJDi6yda
Z8O8RBX8hWOVZQlVsV/zBwJDGIeNqzYGv4YbbwtbajGdO1RtmNvN1F+yA4UaUYmY
wWEkK54oDpAbu2c5qrkeUR1yrjkAFpmbngL1xegrNmpFyQKVMDvlyXZie7CTpbMH
QGyyI4qrJW0CNdLlSp9km8PiGsXk3JanVCFetGlx/nTlIhMzsHHdH3Mk/LklFgkk
ti4G3s3XZaC1QeL4IAFz6smOlCD1yZ5V+ATHXThMVUxcMSEmdvIIymxlz6/1c8WL
uYmLTJoA7nyjvErd1epxkbTbwWj13VXiCn7mzM3BVvNFB+Fzh73ruIXV0J/d4XmF
prkbSXD1UAgKOSBHC5vGTifb2dUk4YW9IqnBtCiIWScsbMFD1AOXge9fxZM7lZsx
YlJXarQXoymElXmTaEmBMnJSB5HHn289M7Tys/VAulHdMm+wi2QNuEvODlAbIbDS
G2eghitL3M2UpLpMUPC9FkMrtUadtTuFGUHm3rwLYUCfQWl2kwU677I59B5JPUDO
BsHk11/se7bPAe7z/+whsHZ5Z3BYSAAkE/jdhCF4SsviURj472kqafNxUGwY71hB
4ZdcJiW8HO43mhiTAkmVfA30CnFvyV4QxQ86Xn5a0vLCmdXTzi85zmuZ9FZG9e0M
bRYsYWX6lBVffFycgu6cMD7S4pEaR3PrqMPk3d2FhVN5+2NHzogEU8VEX/wtL6Iu
2yNlzy/47NVLXxDd5cLhu4jiJsdR8g27nsl/YCtJbugnC4u4fR40kii9o5NAFJq3
80uIlQAePoQ3S9chrazL76Zvzr1fuL3oM2GCgqNmVplSycrXfsPyHgXugcY+P991
kQnqvPkpCgf/xiH4b5feNkmC/7SihhnLD8MctyMjQpR0TaL4KP+B3z6OWkB9Ev5w
Z1npStPGRG7v4JzG6JgK/oeeiItomGoUBj3aCpVc9GGInx5hp5rcG+tAdzGMLUdk
6JJhLG9nDi6SdJfpCSUABxhTPd+C3iAV4xNl89bTw7jRu+VyVRytJlCroDZY4pFD
Bl3PzWTS+kuTUCJXQO7pSnYpR4kx/DBVyBM1FGTNUZvmqQCCxunIeyiiFedkzpfY
rBoCP4EZcEjvVuH7s5cx7UNGcxVBYkNZL46MpOpNsPBVU97SYK615lI1Tj6YxHsK
bglVJE/YwJs5pocjOhGUi9wzgQPLYmkQSEXqEvLO+ZVaCv9Oz0vtUUKeOzrtbPZU
sS1qkDf4May2rf0dLiwiMe9kyNn0Tr9EAaEvynH0iuEM4z8LDA9Wozuu00jn3wPz
is5mW8455czjFP8o0EaRdPNGmx/3+X6/HzICPvwbVGTubrwf1PHrRabCQGa7NKiN
ViLnAqtMde777Jmm+aK9+b0k+j5Igdv2idWBFNyKyIewomQNguINAViML0f7ap6i
kdPqFvkwBsXc5vY4dVupe4vwcssJRSDKL1V16JAr/CuzgRiofVAt9vGz6RtO7iPd
EA3mUBeGNVVjlc1j0Y1Si2AYqQOVWgSzdsJz3vWnIyFOVwot0puoFpDgtQRKOG1e
KhsW1rKJYYQ9EwxG/yJSItDZmm66gXw0dF4Q3lpTg5ALFLVCryEZe8rTmAofdhOI
pHQ2JVJFI9OxUCNNnwTy55Uu8H+qzOG32qC5OUd73GNDcc9IudX8Tv5xcRCt+pRt
a1K2SIqoH2lCbBHRoWjqdAaCrCCrYc7wS+2V97JfB5wogZg0rQ4ULrdiRZun5knn
AEOP6Kkwnuaa995IKEo4qCLLgIiuXwlTtijkmljZzVXp6GkinKwYjejsqtw06PgB
cvv+wDd/QRLWVM7Czv2z/51zMU7zuSIBakIKhmzHZcQNCkkMs65R+Cy47bVh8GOc
WMtEhk6m7mZwl+aoRg6/uqHTqov6jBCytqlCQXmS9+MIKnFADmbyLMDDcoR5i/CB
8Dir6LLkrdrfGTErlOf0WZOy6+7uZooYw1VyyY9ui78Rrq0GZmRBKiF5T2LeLoMc
kOm2kGm43yrSDZ7IHyqmFSza3eOyEOpfVlybAqHKG9aAQM4eJlCtmVptsURfYfWO
VuRT3B13amLH6vCbB+rA9sHzZ3jQW1pA8LzCqvP7TqWJS//e8gnGj/W9BQ4o/V1E
lv8xMp+T3laAUf5sFA7P4t9BFVN61xYInckY1MrEZ5y+hKkK47xBs9gTEKtlW9zY
6QotNY7fLKnPAxGQJtQafuYhbM4zPEy9VnsX1ZkjiqOJSRBV+4dq6+onxDIl/pgI
AyBg3Tf380lX93kdyLfS8ff1oYSYS4D8eXZME5cnB1InWv2VEd9juqlgA/sGh5bg
5r2ucf47D6rkkB7TwS7f0fG7HhVu2gDqTinXpN57QkXYZEuR78DRqMyZF89gNoj9
k4XX4l2OlW6QuW+YXBLvVNR4TZK50r8AOOGGTRVo+B7cgZC5oCucecw6IjNm/G0k
DDpVxisdRdRduvalhCmGQh2ldrApFUNQbnUyq6sd2J8aG8zXfAtxjHmSdbizxoJW
nTQ/iT0fOY1p+EVEqERDEbj+QrGMUqq1vUUiUjIGTTPvJaXSNOGA421P1ZiildyZ
j2lGjjxiqILEuOoOacG52Sl/h7/+04TUoPp+fZN1DZKNtSjXXrj05svWGmpOGujH
Sv47Xst+uf0XdlcRaf5ZnLZr2BG9g4Q9mROJB0hqz74EIwnn9gBnRaIqYmOPazPM
/SI6orH/Nm8kB7r1Svg0LSA+hTq8Mg+Q7prUVX/7JqRYeKFK/XFf7xzy6y//BRDC
YhOmo51EA+9eoPqz6yyve+oi/HQWQpKVQo3Twiz+WgjQmeeELfisI6yuAQGfjptW
6OAZWHSmZsYczs1rrmf7Ch70zEGdtECE5ZonZcSIw6q8MkGVwxOufR1ysKR8RCfi
wguayNGCGi3azCxgnJb9kQ6QjJ0+IqcdF1fZ3zokxP7xSWGIUCWNbA2rtYU8UOCR
1GffioMpWJnv+jmbFxhht2RIXOXBd61avAjBi1yZargR/VDW3aHxJpQHQHf6aCd7
M2gDM7dWI5GqpS+aWvQbWJywSPu3s22es8PrvT9VIxj3VoZkNJ5Ui/f/K8J03zwW
Vj7CgfYkFhn1HVvjEI2NV8s758rlw74+glV3ES7uqCfYUxLKgB4iZM+abMS2oTB4
r+IUaAvyuK92C+YHRxEYvf6/G4gtexIsnadhv50bgXK7IbPckDJwckFLqSuACJhH
X+AR18JV8sjC4yYzbF+sfeU0uwb2wf4oLTem/UpOrviiecHj0yG7meG8M+qKjAwp
5VkntSsG+3lz5ZdTpY/aZJnMw+CMCzmCx/rYb0j//WtdmGKjCgiGvKr3+MTLTtXF
O4ljSaBbYsO+LbovwoHYWIWOls1lvavXiEhsy6GQZ0McSzdeO2Of6o68FwnRaK0+
5BrGmVKEmEqdxSvtvIrnx+IMCQMbyHae+fEgqUAr1RFXYtZLcLLnItzCANVgXdpe
QEH4UhBj/f8hwBRtqboaOeZaVmhrrzESbHbdImi5y9VES4OIDjGmuz8cyjgLpkuc
PJ8CnGitxCMe4eqR3CxAH0QNQ707oydiQ0dJddKN6SjrEaNstY7Ga7yj5m89oiYp
QHM7i1K8QaMDNjX/eWX53QvaJ1a+OW2d5DprBHV+9zU/Y3oKUhTp2qgoPZm/drDD
4l1jodNLB0HFwayNjYoCvA1snVkR89mt5PLjxdM5xy0BoeDvr4tdxDhB655ZzNHt
EDfmxcl6EyFGNat8p2iunPFQorSyzLyWnH5UEQhNNJpNEZZjDZQvPnbq9jOAMR2T
XjNDqPCGg6Zu2HXmh+FY/AJuJLvS5UxL+MbSttfHxYJ9XWfVsLhPhz6IOejBdGov
Qy0XxFFrV3R6THFTExWvPc/W+mDVhtGfBd45vmWLwg8vKFaU47MNvnIqA8nvZe/T
w7oytetzMetgkgXbmVua5LlMv6Yo3xkTiIjHG+ZaTO84S1ESKruXUTLiDhD/MycM
+zHBtkyZ7yjVl/pSpZ62oMVYBGJu3R3uWdBqYFIF8ohb6gqe3xZmYPymaZQ6UfYB
fkHHtreRXs7xXmUN5NePGSMtPRgGUQfM3lPKceuUEZQWo1RCUEg+B0lIQ086K0kI
Qn5vKXK3QZorkCw86oKDVCQGVTO2m9KJQi+YsFtollH3D9/D/dOZu771e1WmIgWb
tDdtlKJnxUpHE/2j8PTg7zokMMhzibaY4nrn1k8tQrkTgBpZaiB1kew5NkFlgodn
CTUkkglK8qt6JEc7PfFmK4RSzXe4+hgO82SPLXyt0qKtRqWhUmX407jPJDDYsSFq
VrBjJgENv9PwIZOq2pDCfPNDUkGBdAQW1i6l3lFNhPu7mH6ULTji9Nx82A49GLJO
STwXU4JzH5K7dERq4W46J3KWyZGwB+r8+nyuFn3RhcAWXkT6pyXmhiHTMKkVm9jO
nUtK6ITEKzdWos1F0t4VOyK/OGzYYier7bL5AGyGthbAUDHA9k/qmi8JkuEzOCPp
m0h2Ynn7BLQrF6azHFdIPnAfoIg8A3y5hDy78WJXSo9Sulh6PFefU8IczDE0mash
vHhEm8tGAdHTSnqAEjRK5A0TgzPf3HazQjNJv2JHAbpZwtLGIazv0IzdvZ2bnkcM
3Oov0rGDYN9ACOZrOSV0JrYKJAcz80chcq6rLs8OAYc8UK+XN3AofgQsF3qylUSx
KTgRDCF/6HV7sRhvOTU32uYqKLPB4L6MXE2vBxT1RshEpBCI1oUEvrXYdlY8fOfb
N7p94EutG3f5v5HnnCJcuoKlU9OTx4WJMl46b9uTF/r2vV+5VggQH8eEAHDmO26c
P+1vdIcVFIl+fU0nERezYzQ2XkZmJQse+OmkeiOcU5jWfA3oMyrucFEa7M0OioBi
djpJ5FAd2NqV9iuJWA47JzVD9WfUzQ0DQ9sOccjzRL0jsc67ZgsONz4JtM3DahSR
hFuaW+0WEbYDnfKvanP0iJHvsvEvMF5TmSi6NXGZ878M+WhXhIzWxPgwhwSMY1kN
YVy4VU+QRmsKdrJyQc80zET6SwiPd0Fkz2SzBi3OG8O/VAPnIPYMXZn3/5UuV8eN
7V8qjNBlwJpwYJV1iw4Mudocj57edvm+1SJOPLPcDa/gmIHmbYYpPrCDsJevZ118
wpfOMxMoBzXwYS0DPvW5CHuesjPkPCp0p3LsDbwSVU9yIp3MOKClVPS0FHb37XOE
hfLxVtc7pzQqbZQl2Z1VNayXfp482PbUuegS77jPDqJ6mPu8FNCq+cuaL8Ray6OW
J+Dxxf5yqFN+xGjdvGnqo21hwiyx3oEf2bpgaxPtW7Ug4KDPT5BUQhn7TMC/C46h
hWJHuPT24hpRRR30s6k8oybrEbDrw5P5QDwiAB8GHNTLlBapLB5kzTwuxS1i16cN
oqOPKMinLaFy6mkkfaT04u8oc8PLuhgOIXMgHePNseWVEKyy5MnZtt5bfwGgKkw7
zBxAkc49n22yJyA6+wNpcCPBPD4b3NZbbT7ao+eSn0J3Lvr2qyd89MSWWpQglAue
6kKteRaNBXIJ6G4zEGs8RnfD3DMbbmTflklm6fDBXOf5WQcRuHLfsJyWzv7UTpmX
vKPsa+2stJorbs+tM1spbBoclL/MWDqiYZXACkb35yQ91QGyFtkbcdBQZ4DRp8od
eCm1uTSlCN0H9kCwjkJY4Uht+S/TlqeWJZerJqBpn8pts0aLB4nhR/XD2lYjPJ5H
5622ftg2iMl7EkaswZ8DF7JfTOI6iD3qbXWpgEQCdgTZ9QCobZ/p0HnnKKn/9l0f
Amaz6xTuv+UPAVPKD07fvXcwlwXYp9BbrVqPQ0OJ4B2iTPrRBRNnTKoy+KTmqtd9
1Z/mkxtXaA3radQ8Ha9DeA4o7h/DKwqpWpQkeSmRkF2TNCUxNkepjYsGMWEcA00L
NxhTOUa8lKrFNQp5xio8a4QdWUFg+irBKt9COqM9ExOZ2WChheGkYEhHwhbeVrC2
fhj24vM8OwTidboRBYVO9lVIlaxkqpIH6OjP2v083N+hDnJm1Nlkl8lViEOIQgFo
VuNYCmFD+UlwAeeX0XPAkc2uhvWVCkSdegvDw2gWcqqOaN62Lyq3pifmnEyWrCnq
RrEQpRsApAZxPMiIIS+6Y4ryAJvj1M1vrOflcbKl0Pa0l4KgMFkTL8AarDRuSNCr
vkR6Yev0gkJLBqvEBUrYDpUlZsiaV34k5LEZ6igqwUHHtNLKXW3nVieEVDQARZee
PnMvxsOQMsuA6XrPrv6FoQ7dhsbhsq69vJwPFkxqlBYYODVk46d7YY795EsKZEp4
cCIHn/u+rxD72p4DrrvLWf6uFfyMicabV/QEbj/aA/tt/EhMkbMuJar9NlUyDa2I
mnAVAxr94hgy9DpcI63IFHiue71qXtwQ5respcKzBbqXndL3RE8H1p2PhgmikV3i
ZrqP0g0LJ/WgeQvXOXIG50w8qG6G6DXESbkBzWtzl2Wj+cugSDS087eAaIO0/+4t
tC6Q0kt6vql3iJbK3a+KrGxlbGTkfVWaxfnsHCBS0akFCar2gkIaZbmYHDkvwKar
zO/T8Dd//9NH16bvF/g/5VlyWI0MKldL+st+grFzEG6X8YkxRnC285RhZ2hTN9cA
rk4p52LV+mK+9tAdAtAx2udBWHJJ91kRzlgfzRE1QL+31C5px40modvqjeHrOMqm
AAu88YmG6hrdkPm8XDwxYx9m1bQSjSsEK8Ov0ILHjWqPzCc9gzcJTT1sFpwPZEIu
xpJYAPRlmmUmmz7jwwiw73CFdrscpU+nVIFdlJ0y0DkADRTu99jmVRDjO2VgSEWK
/yLWty3JvaNr7bvIBAOMoNa9+V1bKjqWZH3TV9PTyj5yabFYZeLhl8L3CipQaROg
KNP7LDIAG8G3hktrW7v1P1OBYwuFAkNbwZRHr3ss3l9s7ExI2SubiEGYZDeJhemv
v4o+JT26IUZJ7PQjNvjiK/pr63DdyZfX1rL+CzjHiPShY70bvWISzguOHTx+/+xl
tN7Gt+ZbSjb9B2rWqbuurRXqQooSjZ+kxZrwHavIMM8vs0D/8Ye+et6HxL5p2yLW
PhoFfPEfNsUqTEVkRBHOOxGUjChBlzPwy0fGarhLvHVB6cwjXzw9KDu6YwLVYC4D
R28Qkh2t7L7/8j2EeoHDF3IpFBy4hA51l8/I6YLdpiqmYVak0f1q9Uo5g7AMZBi4
cTJG844C9cRl0+dBDGVISz619T+322yti9CUastqxcR0qq54/o5NYsbrN7qwY59l
giJQGIdUTjkWEiCtYWHrICKbdH0wS1VkiOUwSiBM+V5nyt9X/EiBcHIbW/fc6qbW
Oti/dwSs7qt9KKT9SIx1J7RSV9ruU6YnoW8FjS5VoxuXy9Wd0jKMZe3sbvIkN76L
uXX5MCkAkc3yZ28AoS1wSb7AHv6Q7O9qFoVwqhExTCt+sm4rU99vPj4kax4DAsSe
em6xlrQKWB5srW583VBzmhxMIyrmQvp1ptpK51/o6sP20jmdK1nSfrf0irNlCC1Q
RCt0ShvmqGKiRwg5W7qqE/pToiPAMrtzEIGgrjnV3ZO6yfBUUzqDnWBZLf/DKhKV
i3QLiWgRaKCjd8i2tsADNAPNIXJuAI0UKEoBArZFrMbtCIqPG0TmOVhar29qv8/g
fne0K7nfhs5f58fG8IzizJBr8sxejQkZaH8Q18Y5iU/4aBvSS94Vflpb+cfH5crt
ny6qAuq8KJP45rUlqu3lGlVqYz59cjIcDVbwcGXqjKQWEpo0VaPjDX4U8JE7sUM5
k912/Y8sIU0piV/mArRPAMUuJvPEfMu3ZMipiR3qZFa3bEr8QgsIHTaa/g0+o6zi
9pmCwHg2xwvm0gf8M2Hll72RvlAKRsMB4cNZqLhntXYfnTqRniZu0yq05eWV8bRT
ffHyvV8SRQ9JRousMuC51uEkb2pygeHzN/K5ef9fLlkXgPu5atT1xRkTucnpEjjJ
2d/zw12PK99NFCNCAzqYRp4x8v1ZyPpShlOJNHEKTB+X/kQlCtu3ihur1IqFrM0n
kcFBuLb0iNCtiY4yYzzHz2ENnwxs6IXT6R0j29w6qaDPaMHNJPzdiXwYpVN/8vWN
i/bVzZkiuUcFOJaq2wXxV+BQ4sTCHcefEng/YuD9i+eT8f68e3keu2YUFD87KIT7
HRf1p2VBu7H+yVU/RQmJjzoI9raXBXFM6z7JdXIR9DgsOcP3xGfWfYKeBQsag0hF
eyqrDUIUSZmvbry7tTHArOA/FV1pRAWk5V2zJ5MSmu9KM3uWpL+fEFNzT+VtdyFH
K8ZMjFuTv9eTcZjKQXsGZAq3bNN9TdMHWIsMlc1KWTV5/8wFHGPRbDGIKMleSBWk
ZNCnf5V2+q/pCpv/AaFJ7WZya+RQw/0IUwuKi5N0bsPy/7FuEEePbgu4TwNxUQz2
hBb1gSuyYS69sqratck4Z6wI4oCQCZm6Mc3AKpu2TSqipmDLDBb7/lM5+LD8HVMU
Lym8oWa5+xl2jOuL/UN1kbse5nboCoBWgBAu3kXhnPAxFYHzFBZh2bj6ra5P+er0
rPpktgX48wGNDIeNHZB/xIxrFYohS7obBmoS5WH2zDMiLhKQxM5Mn68twPU/IKoJ
DA5XObYpwZZPsiNh3SUTwZctNSl7RPJrH1oawTHz8exokJDXxa61Lt7EtZUFKyQS
s/QOM8aYn0rBOQhEaAJPC7aOXJj8RMkKEFHk79DV9bGMSrQSOA0kHCG/k+nhEJ8+
RocrfBiiFdQZj2BZ+etxItqhtt9utIh7aRBytnbG5wAFj0jGj5Xufo7ht1qu6NXr
FI89C1ifHMwxg/BcFqAyFUtJUxKPD/s/fv58/W/HSc57bmYC2sNpzjeASmZDxc8N
By4/RY5GiMGDi6D7eNDtfJQeO8oZd+tpgDGVpSzzvhQEWaRVRlSvWBcfcSnaYNsj
NiQJk9wMhCdG7xX/agel/jcw35+b1yWfM5ZPhpcDEajCgCNytaqvNpFlGEvhMtUF
Tz60aJ4OxlCb+XPN3EA3twE7K+R72neC50MiL5WlGD1+EpKpqAoTr6eLxVvVz1YJ
Ma97tXFYSVOSd6F5kM63YcakHppGsk+hRmvwZyvQthamSVQsowzOAB0CGlPc3WyJ
e0LlwCkg3v8i+N5zscGsyu444FW7u0XHfKUUwFxOVKc2IvXw2Sj9Ryz+4T+I2kIb
NgVCcqOT8TXUl9iLEEN6JBFqXSR8MDL1//1YHroljWpESZOLba2OO87bddTXcQJv
Egq1c8eMSS2XG6snWHieflKzkxI8KhYnkHRexxCDoRLOrHe6zRoWeDUyxQeT9uJO
lbGvivUCLNz+ygW/UjJh9a1LBRd6ndW/tg/b94KlDbisnfUVnvHggFXBWwo2wYcu
03CcyjY5jNYsj5qJRNvFjxXDSyIwoaQ28OBRSCyzm7wsnoRuIh36wzoZNPNLSH0K
fETMo9V84AwABSg9Avm0pcNJan9VzgzMfrDV6FtKP/mo3KfjXRJn7hkWOoO3xKmr
DUJoGHQKpCO1xPsSnfcYTtSDwfGtMvuP99sgj4PuJ0ivmOvdveXUvrfneRlNiJAV
q+RJdOfVCjjiJMdXZUPw6yfMK2jw9QUF4g7qPnVmhiqDvyaVDUk40N9WJcID29mf
24woI6Xu8k4X6w5yuYucPpETXK/101UY0j7BF9wBqya2mnqK9xB6wiYbnHIc1IXx
Gmd3tA3unpIiuhRSgbd1VL/9CgyTHCKeJWpoBT5FP/p9gDzY56OV8/y9N/a3GwYM
gcDvH25I97ndDecP5NrDO9XV6+oG9p/+2Z6rFhANx8Ydi+puqWH82m8sfRkmPXSp
IGvApI4yFy+Yve4IxPo0/I/TYbU0BTCkVxJvvccjwHOk7LEUCFQJg3WrQN86Xt8M
0hQACpBIdC8FaM8Xu/W4C9Wu2705BWIaq2OcLvR8oYAr4EByx3AQ3BUYgHSdCFIh
AlfqiyYhpKmKF0KDpmNyKODmqEsLYBjATbEZNs4QT0Px2waymh4DnsQ3LxR23JQx
5SDTueleLuAUA2u7RF8pFz5mRWU1XEy9v+eK5kfId97VohmXrEZwqvlIEjfa7rlF
TPvLUAQaxZDFkodY78bs8MBb6albHrhWX0nf/Z/gNqhk8+anGrLoAjTY0VL4jg9B
0MoRcLDF0KW9cEzpoX37hIpv/qzUmJbuj+TT0LBjY39vwqGTE5I6iSGJOEmBES3D
R5yXZHdXK3WIQrJyoxZG0kQAjn2gBDHET6ifPJpd6y3sLqGw6h/1ICRRqusePHY+
IRw7+vE++Elbv2DCFHR/8huwf/PGRBjjUE1J8tFxtDZXr1c+p8vr76zcaJX29IOm
xrc8OJD94M01W1b0vgcIfCoK5bXWON2R2ExfXFKPK8F4ievnhxaFrPClg8ObIbUX
AnjljU04c4dwlnZxGojvGT6l7+lBK6GhKt3YH4e3ouuKBBVfLfEGtMwK+Kw8HIm2
qfCgQ75oVnGlP307CvxRJ3DpialMvAIglJmj1c6+eyyfbEEtgF4r/upUWbrov4Lw
UPAQubXmLC6cJdvbVjtDeobsDVaZMmIJU0WJfXpRTH3WrhEJAKJmcoX3bquMvlij
ijR5rckFvGtnb2O52zp2W45xutaRd03fLvi2B5mmShVn8gq+mIals0cUJzAmROgQ
zrc4Vs/EBs1ZhvEWD/axNPhx4iiee/3xyxelB8qG16Uh7/Roybzq6xbq2bSM9ycG
D8jNqtWn7xSk2QFFOznrQeOF6/vyXp7gf5eaCMgdNf2kX03cVvw/zY19czeyoV1S
AEI/GTO60P/Tf+tm0cv+4Y/OM8HJhncZPDQHeizPVETGVPtiglptsEzYd5MhcDzY
Jndwt5xmuYS4isiWsilIYbZpo+My4u5TFCOwxVypai8Fjzmpy3+0fykTurIdVGdB
0cZfwXKiQuubp7iYg37gxX7pkkx2kFSk1vIdBqsng9VCLbEt42nD6JchQ4X1sOsW
5b5thoDoCh7YZVwKWj+xyVdLSYDZuIcjZL/aMVbGDVOJII6NnUMX4/rf/BDRsAq0
Ox5N2ChxjBDAzNcfIPgRmd9zKUi4kELgjDNictE0Qzw+6JvHuFMYAWnKEfR+2viG
DnYAoAX+VTG5EEXxu4WgyUP2fRG4TPpke08Mc9iDpRLx49U4wvDa2l8o7dAIcQMz
VcTFzLB0Ga6lDZT2vCfi866JgtqtizLgA4CMKuGSPfYX7yUzLXkBUEmxWi3NTqnL
vrw6Oy2GYUdQu0v70xWJ+IqhvAvNTX+Pn/kf4QZ9lsVcEQYbORSSDq6U5XCML2FC
mY8LB7B+7Hpd8bB2XVu62shnfVDenyig8Gr5VZhhsI3VYvtHOFZjEkzQ7gwQnJ5a
PErupct+FELmDNNA7+h9cuT0YOO1yF9bXXO1cwB3yzOmSOVa514KPb8t+TaYZZVk
gLXN6sqGErRZKmsZKzjCKbRifyXFhOcCotV39OJnI3sgQrrF9zb1rO6MnzXdLRcD
PxXaiQTi4cw9GyoTW9TCx1MHy+dCCIJOo3LEq0WIWa2aAcJRAcE8SN0cxYBO77sj
rfhjdLSzp4AiYs1AQpQIMRqLaUvRXPs1iFYtp1WbXewvR+4MZN6w3omDjmWDpQvX
QkV7M9rJ1Cd2qAYGhq4Qb9a0DiThd1v4pDXloQKDATYnV9x6Mc6KUSFaQPq+VHBB
hoLHuoXt8D+m9jAoHcohIKl3sQSE62qHQdzgL4NC8op5RdwcBRcOhH5vdcfcgfGG
SC+95YH/bsa6OwbjHz9Wb/bxFJLw+BN/iUZAqN6vZDF2l+QbCt1KUe4BtGGvClog
tjYpRgIF+Y+HGwaUARJENcN3VfR7pkKko43WKxjPcMZ7/vfm8kIHshfWepzxTszc
AH9trV+LqhO7miR7mTcQW5oZJaTbkchWUFMfG3gk5qnMOevPzsSoxvdXR6KwSqM7
GOj6Ewa9LUf/7/VInbNdDn+qvbC0yVcO9Z9DW4ebuI67SVPEoEf0gX+5krwkw1K9
ZVuQmmjXvUUZsb0Yr7yPnh+z6VX+iQMMZBvUUbb1qjBrCbsvy+jtaAkYfEiaqvFI
MCpzoEAUAwJd3MXLZte0JauSvcWUJrfXmtho/D/vaNDXTGlxdxe3sra1TwrgFE8f
XrQhI0lkClEQ9ZLWQ4ebqGD8bwwy1vd6kHJsTJVZCSW+DVTi9E3LxQbeUUit8h9b
tu6dLgsykxKAG1anieC0wto0I0s39RTUS2IZ0nQ/E66awQoF7pG6hvs0LQZ6w7fN
Tq+NLNkgleB4X5UQtcCpV1tQ40YIMocNG3ix2VU3E0ZKCMN+vxANHfOzgOPByStG
k7E0MBzTFdpbzyBfWFaJwrMduy+D6Xhu/FrIDPJCKyCWElZp8NgKEU3sSXIHe5Pp
JPtM5M5vyoykqQlRSdNx22gc1tOvt03UNmAOULhmEupcET0YmAfrVymg/hXaL/UT
YA0rDsCu5WeOnBJGWKOj7/efLic3Hk7k9ZmCuSK0rBwanXypvIplCwaeFjTwCR2+
Za5hJN2buExm4Qe6apXvk+XrYoX0n7YSF+JjTOAbNOtPPybD/FV7tr98xL93RzaX
wjDz6EDZo6ccdu70FSl9GE9ALuEvLh9J3voPCQeytvwvNtpagnq8EoYv1HVrz1+Y
cuKywN5+6YjsUzTmHJkSbJJHspVP0FxbGfhp6DrAsfdwO8OYlDxHBwYCc/Y7hNi/
kb/SeSTKVOCRIWVApCHRIpH0UMsrwB3kW4qV8WqpGUGx9PtwJIhW/IoJH4j5YlP6
rqMKdX7vconn1kW4lZeFs0nBFJ9/GykD/k0sBO981v24tZEjjLQVjvxeR218tx2d
0t2SMImD31Rb52xGLZs3kz2Ec0iS1FUqVa/HQmO4q7U4HdJrIlpg9MhPbXuhq+WF
5z5YdZ1VhSpmnChnhC9dJGN91OTWTdWhIEa8AhDXeJC4oYN1FU3yNaNO1241yExt
BKtL4i9NPgbRbBrIFf+vreQefGUjLp0dq0h+aj4hVZT4XlhiXXx/rSUrgFvoBjSP
9yhLsP9HplWfFC87hpAi6OP+RdwiSrPCus/g4v9eh65IyrG2B3y7Hy7e4mMxss5J
OL1G9q5V5JeXDCNjG5dfpVuO2vI8mo+6FmEhSDOR40ZUEPJOPIcLS0fN845ngro1
SEzqRDVGA+Pl2FR2qEkeF/HdgOZttKlliu642SYUJycajDFmV5Mr7elB94kFFp+k
PfHv/jGL6qE7RSaJO6h1SqMD7yvebGb8cMi/vZSyxH+jwz+Z1mWf/cfEgIfA42eS
Hzy9BqstvI0lY+Ig4XWm6FhzOHEjcGoTLjn8cwsRBqgygLxr8C4ITe8odQHVeMph
B7fFRVhR5+xHI2bCKPV26J/3Cr3/cYQXRoegBgcr7gdmo5FK3kmWFDz0X05On52n
FOC9GV423nt0H/B8QgbJoNdOlqqOTNExbwTEIwihOnahXW+wp6yH6A7SjLqmn2Gp
vugZ+gm14pASvUisYUDtvhi8a642iOVPLM81KnnDyvYXv1RB6PUr3NOF77PIq6iT
1YBMQJVFLnx3wGGHud7OhTbKU8AUHga/eC8IjEomarfHzF7UkNEBJj6qYwdl1/wN
WI+RHlIpzwsgvseImxYhrkP56b7imCGCSV372WKXBrwQkpzmkI45JGVARzVG+F1B
m84wOs38QTntYuyyMZCi8f7Ad0EB0icxBRnAhG3GP+wdpDiz6famktGm7VnjSxTI
gkEyAHy4NmENarcDNMGLDl7albwbVhQ/r4Fosw4iUfUDV4kAYVDtU7Be9LmrPN0I
YEtSUNvl3fH6XLXOUjjVXQfZQEyIvAu5cwHvvn0DIjfUosNB7hwVHg9PCYOnXTC7
TKaTwpi43AbAIHZ5VuLhSajdcn0VbcxHJTFv1ysG6mxdWJ98yIda6l0R/wYkcsJ3
yXqZdIvgIv1nNVgHULm4SpRH5KbheIHBTXkHuufjjy0bEONQ3YDygv8eVysFh9i6
gQdhi0nuQ79LNXWd9OurO/ynbmNgFXxVoMb9hbeBlGVzCV3pdd7Cz2n9CEsn6pl5
rX+Hgg4Ty8bgvlQiDHP5EElMaUu7M3gPLLGfqnOcVHjvbaYDlwyVr6/JAQEdpxvk
ewIIXuC0REk4wvPPygIGYGV0AlsA16SYXwqVeSQsq+9TxEtJAIFnXHBAW1kAXgIT
u4BJvImVqAmojeRnx3w8Nh+WEyKaUrxsCoNJp7n/so8/QCeWCahiyC5eVWKv468q
4ErRlh8j7Z0JdSPfUzKE9CAT2naNp9/5Nto0F8/qvIOL38pfb0MLR6MLWCiWgp6F
Pq6GcI4GFF6tLUuBugaauoapcDryBgC6+0bAQQLykiXCr27FZGJXyRfaJ/cMVhy9
psjiOFxFAIe7QW+oUOIVjm38U1251brh+2dflGGmwA6afF7xSoSH1OcAC3FWQuy/
uhu6B0HzOpXE+pbbi8W/uUxHMvnRXNxT2ly2RHwLBOTm7O0qI9gb+yfNqWA5VOfx
k2TXfOJDSfhWYEyLTshlA4RPKP09iB2nXdnIG0olS/I1ZMZEfGIIpFqVXW1QJdlQ
yQYXQQY3DISkR5EbBaabV7jNDXFucR+X9AFJedCQEJKSrCbkt2pUok5IlTnoRWvK
JotNHggRAfBsakcGSp0TL8Vg+lr3nJj+nOzFr0L7VLeMuLPulRcg7/+9SxzwylhT
NFbXZ3FdIb6KRolK6pW1R/ld1Ko61/y01fNRdrHNbBFYgOsnqP70InlGAL9Z4LMc
f8zL62obtAz8uVUgYUJgaz0vt69vp0rrNPsOmF7iBF/lxpSUIgKWRLSxpvLgYvfT
fMv4lQhOFQsGHPL5eV0aFJdDWsBhcGaacl80V5/lhSRDnf3rFafPEriVOsev5Jyu
ULwL2z2k337eiIPQ53XoydwFvoJYPp1i2BXu5MatlJneon6AJO9HsRC6Ch3tg7lQ
GKgtFdaerzs9VX/XeAZckmUfZ0Er+j2sK+f71K11AlN73MmCnU1OihdQII83pZAD
B4fTky1WUKT3nkiZetoOF5f7aOquuyAV6InDHT5l347u1ZYS9xn4UXqyI3LT7m05
iiDhGsUZ+AhU/jAqhkDwddLADn22W2tCAZfcDlHbFrOu7azMR5zDIqN6f89CX9PU
yBSK5dAjkJsjPNmu7Tryr0TC8S3T+pcf1dmphlXd1buSi31wbh05ZwNsfRurj4d0
nheddOePzVUYbCb/TnTGkntjyz7LV/eabg4PmpbQOp5zay1V+a26VUzok/deIBHL
4CYRYbzPoNwpEwsWynPJ4+ZsQcBpFAM+tBQSeIZGbbDZHHTj9T9b07U5mT4o6Etq
NMj10rtxNl2Ip92R8aFkEPIsZ/NjnL4CmgfxkpHJJvlprIqemDcYfTxp2SXdNL02
fXoAOWg/j1ZqqGgL4OR56Q1nUfGGyMLGRFhORqL3y6nepM1ZJSgWRw/A2Mp58Xrx
8qnF2RQGQPGMUKJVh9A8OEZmdp7Orxt+HlwF7a6OBllbHDnvmnVI3HS6HVjXrqal
vUq9ncC9em/U1nQ6quUcc4wOhGS93qIXOxl9/YG7LJgCYuxmLUXdA/ZCynakGMtN
StlFe4wUJgKGDCOItMfQy565/9LtV6m5xIsRpbzfwNwMQK8lUj0Xeif7BOZEZLMk
PlmnnsGH+fZE1Al0DG2B250U/5kcrCsKu8kRbKxLzUooEY/naCFoVEzhHjvrgKnB
AXaus9x7sOHiyOSXlJXq/owtZh8i6g6qqtHKyz3F/Ki6dZiVetjswsU47c23Bn90
5IdkfJMZiawFhZjTL1DHKTiT8+SSZYXXnO9GJmpqhIaUd1q8wcuQIDFuFwJHE1Mw
FL/7SZyiJk1KJ5iGOweKpYMA9QGiysBZWfL1DTh/UrcpVf4Wdx4p7jQgROnPbzk/
K6urEVsqEDvnRtkWK5TA/gmQ232Cv0PXoz9I3bGVDPiCPQHa3apCLA0lMwMvZDio
Es0jTVq+fSn7hgrV+xr/aUuzM4455QOajnUx4NHSqIaX4QUH4lcDsxBWJKAWuCDL
0BqzvgjitLc+evSRivhg0TwSG+jUL/mpnoRGsR9kvp1kX4aci0WY783KuDXvHQu9
XucBjiJgk4yA+qD74GRa8rqdkdHv79Cfu6LnCcTK4dNjRsFVJYwS+JfRt2jSxq2p
3h3pmbJkEBnuB46AAZ1lk/QeLph9shQhN+Jn5uTJ5adJn6MY3arCasB0MsUNHqsJ
IYif9SJLpuM2CfKJS5y4TdD3wcP1DYxQy0DXIFQJAgz6JQvjCPNsYyIjR010RraJ
zHP9sdfONJue5fWJEBtRO4M7mrPXsfmgm180BF4yBiEcWGAG6GQZDmmB1MU0ovx8
EDmlGnFuvCoaEyR/U+q8rluPbaJZSte3S26+mDTKOXjEQIYlnyTf/GCNZF+O1j7G
fDXcRHqXiH2QvWJvM1Bs5aGxhnXRGgmXunmjzpmzMGse5mhMnxJjVpNS5/bMgP1Z
+rrMamV9hUZGI+wMdidjPS4zdpJ8rN+EdAFToSFXsD9z5QPM4dfoOXbeaYTiLoLy
2qkLv7t7Y5maHaeQdgdK6k8ZsXJTrPEDI9KPM4sTtGtyqcEIy7jwU8z842/GJv/B
qk3ZbRipF9pqG/UuL6rQMPO/SqnEpiejItSJHAHSDtzV6foEy8zuh2meBkajbCmD
80x7PYSlI1f9VbTGUyHSTysA04zNmufT/SLQX4cBeRHk/ZO1GLpWm751btuFkPuT
mC17PJy1bWUH9yHu7lDVtFlbuW7JE/kAKJ/e9T+RtV4uCkTR2IuUb4QzswMhUdKj
uJS5HTOjuWEQPHPO8I0NtWDkTexAvAxSKws1s57KiuAzUz6Sn50xqdBKU4QtxfwV
dnPWT8I1LJw9NKIHvRJnyU0IW2hYxn8M2tbyGZES1zUH6PU0njXYW6TiG4yFQKz5
GExMcJ29UyvYlEuJGzCNDQQOEsG/XqbTXq2k5y2bEX6fUbZQ/PGHClHAHeBTI0xi
vh1VDvOwUxUjV78/PcJdmYPE5syppnnvI2TZnzkIKFTvm8ZKbLBboyzR4iDhVbZm
Dkkh15W6M5pigFxelphDGRE4Jjcnej4v0PywuASG8VmvtkTLpFZNqf4MvcbpJDqr
4fHouRyxiVH51+Ca9W+Nl6JMmQRBtWiepROUjzKm8Pj4XDmQa18TWImQBfXylzsk
HmABpVxZDZxMVrq3Hcg4DViEittR5FKxZMAWTtkS4v9LzlKPTEbb/syJX9fCN8/8
Lcsil5uNj74+M8ezaMikJnVcm1WvJVfHlgLj6DIDiGXXIV5leuU7QCs3TSGV7I0L
1f67r6rUcyuqt4wr9IsnNyX462X9tWgSTFR7iGKlzG42bNd75C2gMjcWmAtWlTWn
5ngNopXtO1LHT+2W2WcSFfIltLvItiWB4aCJ2FEHmytQ78L9GG4ZFGb3MxYS2GuP
SbbWZC7+l5i3MAKyj8jt7LoNc0IeD3UXKX6fuPZyccVeutR4V4CFNpoAEw6NbL8C
bCZ7wjox5UqRYzKg5M8miYAVyED0JS6cVy1JAYc5oIAgyWMbn23xKU3qxIgIQk+C
oXUZvNtBW/NuF4y2t6al293Jo9OKKvqd9bo7YgYlyfyilG1Yrss7XcLDJ9kzeSR4
BhWJJ63B1RW1JZtTqHPdKaR2d9qWdBUEOTmpm70M1aWKoTRRzmB9wPGBEh+vy5SU
SCDIF7oZOfflpi3te5+qix9lxFIfUKlkj8+CZjI0OM7rovwCkKz15xnQWhn1L81D
jgRP31fI/MAteGeot9hK5IvNIGj7XJo9COhD1ScgjNtdSM76SErJoltNBLU7h3ad
R4MB7D9U81lbdB/IDbdBfSoD+0ciF0WVKTq4gZyC51qwySgXfSgqxcvrr09xP0PW
k51CWvOE/minJMxjtJ+kFCdOHzM8aL7vlLrSHVryE7oTJjmBGmYfNQ4KFz+/T7pe
VDZU6uuwZpFDRF5NLMpXSOZQamd7uXdOteslIFIO3WQjqnjP+y1NHS9Q6QZtKVHn
KLtqUxDXuivYxMldCxo4O54eUPaMGbrSyk1mYRqA1gC7is5/5gF7+2OJJiPByPit
qdmTXmVDrO+TfrIAtFCk7scwCOTC+hLRU0PaWmE7SLsTn2yRsTrt8XOyhW6nwTOq
L1amSPDjUxUpZyUZtBmPg6/pO2L5DMQNmq4o2aHjeUZe+gInXOE1ViE1G7JB+ruM
PAefBqAnh4IJ3AJHoaLTCVIxLCTUWWGaTVfdm3W85+NYWF/DfJpxvRzz6KsLnVG3
kURQFsxmplneApaOagBELQQZ7wqCPr9fSKq2/p/mwyaclY9w2uu4UOI1SdazUYcg
7x1SUyzZ5TUsNy/qkcWvyiH1sh+oIZaAMt0frTkji7f7kNy0oBamPm6nqkFajh9F
XZeryt37lm82S86uhChylLBCU3g5+ubyBSMiXRzzniLTtJdIUQhKjMvwxJ0e1gvC
J06g9fRuKJM0GtnqobIzRQsSSTYrdTt2yA+hqwiqzpg4idvqqX9t2JHhUuyaCQVX
Ngd8j7S5Y4MCGB6IdV2fx9Ee39pDxV7C3rSc+n2DPadX6XxD0AZZP1hfwlJd/rz4
79mWmrOhkwZuJcyxL103uz0NY1pxPi4F/rMPAxHpQb+mS6FQyTBKSioepMSfm7Q8
AZrBGvfzIPg7T2yy8EAtZXI3R53R5gz3j6GOanFBfP4HgTQdBxjfDMBsWbpJOGy6
aLeBbBjhnYYP/Rc7GxzhEAlKYk6bhZ4rtM8bwNeF/WlysL+x3rgQ45/d32AjLpmN
d+u1dYyVxbSFTANBQNkwnT+c/gTHQeT8eOWUAnzgcbfS4+JWOfERtBW/rZZzBBaH
sZqbibYcPGLQ5ZqMVBbl6VeD6IZTnyoMv53wYIG/+S2Y/5t/Xoo30FA8eg1z4AEt
QFy38a7I5wyPnzGIORsCESGlzEHX0YJXbLXHBtb6bmCb/hJJ1HzkJan8vGJZ19N6
SalPXa9u8FAwsJLHJZWbrEXySgJsPjHcRzda936osa6IlTd2vVrJMnhpQIjwQcgM
GWvoc/QSiApxNAsJFMe+QvRvp4hvFUQo7C5D1psay1ugV5fDYq+ZeqWEdzRlp9B/
Kq9NWJLWsWQvetg8ftE4jVJI/TMNxKYNufuwKNBYs+uUFTHfOT08arris9Lpwm2s
ESb9szfdV2AXaHtCYThMK8A6BNhqZ6CgHmbZWFb22BCwLU+I8fTqSdFFTkyTTYrP
PejfvcauiCsY1vfabogmtD3pe5mBfUUVZoDWyRtBDJxQg4JPYb/dn0rr7mu/HaOw
Vk/WLbAlYKsDpNspfVICuY32p6y56Wwdw73crHgPASgLAW9jRK+b/ebdNSKK//+l
geEqz1pA9tr36DMMXM0PlvjZEWp1im70+pVkHK4obIO5S29fm34p29/Ks1p6SOWd
R3LK6wa8LHvMHXtN0vhGNHI6mnB3kqJrkLtoUgEAADHXPmczMrbag3V71efUknoX
FPe3l+lW+TLZRIiqKcBV/ENEK8yMbaMVkWwGrkKNbu56GJccohAdJazBQ9REcG1e
yGnXXjWmeVRW/4FZAsRViHz5AK0qVAXr5xSHAWNUkFVtB9JizaHKzpRnjFr3Jecg
gvrDFf7mJTpURrLQJWrLTvITn8/jc9ATbA8prM9dj2wdSIwEaodNOXo9x46h2Ms2
Y2s4VVJcsiEQiKYCa3g8sO5XTVeIrUgOw9a50Sv5imyjMU/RYIEs7j/RL+dw1fHG
VDW3VDTyylMvZPa+yj63X1P4ePcH8gZbpsZhKLREWv9KgCk8ZBXRiWH2qzVpMRgB
pUkBnFsHjswVW49ediMAYT1+7ZZky0kUEDqnybrkDnI3Jy13tRivPq9UApoeQz1r
sdyz7Ef/O5n6mfjAUmwKY+U1jLX0+MRVuY2hEJflT/Ub93RuuhMfQMeFgk7hb/7y
sgOi07CZ3nORmCLRbWJf8lRNKNOYz73jKXBXcNRVuSowgLkm7ThvygFPk9ZArw1p
Z2VaPVD+Uvlt6qU2jWjCK8PriO3SiBFQvXwGyMq6A18MQoY6k04M2jfWzFw+OYbl
QDMvVSQoamv2BR5I98oM9iqCPvprHsvBEBZiChk7fBxIiozFOk2RNe350/ftQr6J
1zmFJLGoJNcf464pM83zaxsN/co8/Sd05sUw3MjsZ3YNaTNhCFMGhzDBZIBPE/L9
fkvpFds4t9Ue8vRFGFuPRwoXeLZr3qOliRLKpiwEh+l+SclJ8ENMRKCU4xzlorxo
KwoIlfXhaGZXydGbsLN1bmUhgeAHmb+U+uLIY/j9oXD9neoTY1TPfyzn1sznVa7i
KfV9MZkfjXMjPBLUEW8a5lCH/pXrmzvZFnFITjwOgWi8BwJVdr32n+Bbj45d0N2e
MPMDLL/y3/BwGMTBO6ZQfriIM//gtnwlPBn80Kuior7gTuqZBM5S6tWNkqglwUfq
1HE3RBISFngkc4gbUJ3nkLKbD2KhlsEbZXeLImz5u6osenU3awX5WjppkwtBUTTW
bXzvWFfossCHMwWO5iUGfC/q4g6ns3P3q8tZwo7IoGj+Z+uFKUWJw8/39cNETcwx
yu9beLyFU8cMRv3h67Rj+rUVv5ql8yOUGtGo5DROBkaCF26kmlK5k3wcaB1xEIzw
p2Vbe8sEh0qTYF5G2iFER/IjnGDxRMPUnHtpA7b4G1aO1cUVKVnJLeBwKawcVIPh
QBo06A8QMLjzfZGvAluYAqrg495yy07rGXvAOVTc6PHsRakJmadwue79jVrAjpdC
rAsjHdFUILkET/ulWmiCLOe0izKWpqcxtJrLj9S+FRPXXPJqaZsw6GDBJD5k5db0
0osk1UyKio4UfehPvlCbjCNn+1oUCpj/EyPZhBB87oDxhUbjt3DvL8J8JxAIeqSt
kZFVhMMaMauozKEW76txFVhTIzhO6FmClGLR3A2HDfNZFShJ9MnETTkBfVIo5nMN
ojJhPwNV2+j43kZ9KpNZOSr2CmRVOOEhLuJ9h0pvFOhhIzoXvMARHJMsP3xvvRPa
HRZ5CcbclcG4g1+AiObX30PxBza+Xmp146f2Mz9723I2pVE+GFUiOmV+ffmfUncj
e97cL2pGR5rIV2pAdgdyAUPz9Y448FfkhIxQLaOpaAkc6VWOThEfAnMy5QPr5aYZ
WiDczxWVioObkmrF5RFKoOaNSKRivdPNT9e7BZMkScaw8p1e2AZ5wxWHPJ72hJ13
//RBRSY5tQGGAYLjIAHMdb8kfL+mRbDissJocEH4YjMwuPBoEBckVkh049De8P45
jF3BQchovLsJJOg2VvTr1Q9ohWryhjOvnEZzWTtO8lue8Ma2wurQRa8FUauaIm13
PwkneOn1YJ/JkCnQHzO+pyFHlCBv3xOLpYetphO3Lfe20LWhaAWHSmEPVo6kZ9YB
+TkET5ylLqtSYjnHSm2oo6idCil/10DTMqdNS+hVnk/8A4l+I3v60926tKmS7E3D
Oc7YzxxV+La+R7FY0zy54blaq8em2rUOYfkPWy9Nbi4JOqr78GrQ3EeSGAqUd7Jv
Q+A+QWUiY1cAG2ubgZK5GRIcd5bMouNpfDsq+3Sr8Sv/nEADLnj76iql280B7CUq
jEBsNeHqXGVVzxEqT95g5qHlMgPTBySkLj6a1H51l2KSCedhp0z6eYCU0nvALQg/
/VipypiT2ozNpOtFlHjT+0g/ywIJ4dQjOtphuLmJrKrkQ3UR1xdiUTH0ijWjgPXN
IBJMdubnxcWUHGoKgkLc7+o8MHKQJMcT+PVE0c5qNrzCl/WbvdQjANjlRstqyzTL
6Cmrt3fDwmbhas+WLZUH9mSAGh1c9KWaSIqJitKKTi+3TDmmeIuVDaIBDPT+DqwJ
eYjoKSn3XlvEb5JxmcYRw5fhUmmNW2eMPXB7pnQ0ic3XtV1b7r6OipelW5Bs6DO1
CjTiA6cY238ga1CVjvzEiTjBZ3ko94/ej1wVSso3K4CsTldwqNP7WPottqOkDmdB
acZ8HJJWL5KcwFEdOF84NcVrYRKi7QyaXphVeRGEP5SFpI+xcIdKb81MrrdOVkmv
hMbWEFCizAocWrulT1hUrf7YXS46FzdGa1UEyBqzUFaVCpvQptFaiiFlOQ73egNe
UmhLXp7wiiBX6xvCXRm19NC5g2fVIqSXQkBciYZEOiZ0KiadyuvVWHshq3lXyzaL
8L01Zngy3Oo25Hp0yHfnB6tQ/L7/2Hq+cJMVd8R0rh4LGodh1R0jRumxFqPH2Uvp
fFr8SzYZyO9spVRFkp1cJ59Vx16i8HpeO3gH3c6v9VdklkQrni97h+z844XavsZW
4Smyn3MtlBYDAsGEiHkY1d5p09DizbmZRqN2PYC4nk9brPtX/28tMB8A9IdSy+f8
HD0zuwzmnbXIoWCU6++f/It6EBq3TllMCjHLDJbU7fTxqdR0vpbS/FtARlqsyPLk
khajjh06VLt/raL98hWo1vG+/AC+k8aI960OZiN1HtwVRyjzVkdxlDRhXbOKD2tM
ChRa5giVJSxx8CItASNRRb7ynlTd5JN09KPvHoqlmomL+ySC1WI3XkER17YCQQbY
WzVQ6Vrff5t4lP4TFf0H4NGiAmLdnv9gsf0yzH/A8b8xexV3mVZcpHrrG6sdANN0
wPDJAhI0VA9CsVaJfUIJGXlZ4UgHIJkWPVbuoQIO2AFwYfVKtlzZIY5A1JfvzpsM
mMbbfBFJsB6yiaenQPJlfuWkGFEz2lKLg2UxGpclym+zF+spwXC5sJNfJexvmv8M
eqLw/UKFn+jdResrX5i4Uzv+1Y9Ea4hoeDpwfK3ToQhin3pZmgcz2rq/kzJNhqbx
tYHF891kI6yVEVr5OjjPazv+3QEIhD5PQ6LaLJfKbBosPKVMwW24Rv7Q8cCw4yq/
GSYZ+qvCXvkLC+Y5Fn9URu7lAZRfhZwrf/vlhRgLBZEMlI25Q30JRKL+ofw54bvb
t9JBYZI+T8fuPrmvKn59phaGkFJzQWlCvXqda/xmsF6YxHj117wOtP0rJ47Agq9E
jzyvax6x5B39q3TZpmYx0SMJtww7+n9XiLrCXDErS9w53iPPfd6knKS1c+tWbx2c
d/x+5Bo7avIH2zhGMf430wU+3daJ2uY2N+QBpZN4kSQeXk8iMqL7Jri0R30uqfeT
wtFYnQe7MfcUqu0illxM8O0ST5rLlYjAIQ3/wsLZIJmEAon2scoUYKbov6vzlwJ8
bthBzRGTkz0BUKLfCIDNnLcQsJzBto+lT8DBHz7g3XeXguTe76lquBts8VkzcVwh
sCgbUyVmgaVkK0X4DZIas9AeQQ27lLrTwTKaNgQa4FvK1j9wgjrsCYcZVOJRf3GD
J0qs4vrrJfic6x6Xygagli1HDUDtSsGZ0/DaWJur1H1wZPAYDdXCfR6Mp6d3WceB
SCgBAkwTUedSmydUUylWCzhNITUy97h5HP1cX2glYX2sT9XNLkhm/hvaP3KHQiz0
l80ozcaETOyNoxSKummocP0fctPLqOSAkyHdAoXwb3tXJivUY+EwtptXe7AObzyO
P7nqcxz4/xZz47ijrjgK+OpiDUsaTVVJFXFRt7uwLsCMP7md1m+dwqi2N53MUcuJ
MNvYqmc3sXSy9il67PQK7oyG0Ew5ABBIXuK/oS82IYUTX+iCx6DfCOX1OtdFGKFJ
6fx1ZkxHJpxP2snXS+bBaZldwnqYrlQ+KNoX70/ySB+vVFj6h/6kF85j0IgCSGjI
V1gFf7kGHjlgv/jSOenjM2ZSWIpbB81kYRu4zmOyZQeVn3Mc7a5uNv2IpibdpJ6l
kBJq4WPT46aXIcJMKE/t0NT1xcrw7ztrUMV5nkQuwd1WGOdKCxv/dV7CpFp29PT9
sp7girlgSsQVHwTFNDrqkRP30b8nI1LO4WXzwCjgpjcanWfIL2zBimUbtkN8I/8S
v1y7A85XwqRjyRePUlqKpLbQ++NMn0OQxz80ZKVwrM+yDfmgH7viT7zEprUIEPkl
To8stM+skaHJ29uRRRkhsr0W18ExSmT4lrwHuI0jTb8IdUBv8XM2zUE4EUmSZRYf
2yolX0bOfqB+xOgG1S4AduiBYtNA3dYom+pOYejWlzjSXuzpDn0Lyp0sOmL2aIMp
XiFEGSjmn9vzWF7fpFnuepi8p9pXj1KcZC2MSjn8MTN1LtoOUmjgWboWK403E7AO
s6g5d7vDnnsW1VJPJ/fnRySTVMHmuT2hP8C8UkAhD6QZNch5fv4fxIazjKqjExkN
hBupbjwVbQ9NHvEB+B/t0n3OettIP6tGPPADF/4nmRzd9x8KGOt8xA0jWqBiOM9e
ws6GURXkVZMSMw2UfQYrHJm9nVyVCPhVD1yEvLekiBMS4ctVcqlBpNLXxE77VrwE
9WSwwuQzMdpGbTyselSp6oRO6ImBqGoTNAqjW1McZKsZRTJH8l8HesE5Gsi7GR59
4qAIEFMC5oJq+7w7uSkzPK14vpJ8g3Fm9/jbt/by7jObDsdIq2nGVGT3Yn3d6LYR
IONA5NOcdFn0rs0LIfy7MkhQeF9kScqQCEI24p5apO3/3k3AgqzfD9L64/J1gm5q
nhogpEbbzkBN8Tg6d02ZNBzAWzjKA3VYxdEtDtktaprat8FfCt2oWNZKeBFMjW8c
nMv2HsPSMszwlV0WHBhMpCk6Qi18v20tOQY5pk78iJF3jC6QBf7kr2seTjA+n3lc
x3xLi6F367+Y08WuJ2MXXa2/CEZD3BxLQ8KFxnNB/ygi2dKsF9GAMsGkpn883vIR
RHn4kaS9CMC3pASeldpeQsfwFVFxO0eZulRGzotl3a0AbnsslbbKVkqPhZ20JNNx
PZR4xdyPSnVMarLg4QAN0FqyHJYegD3cGBjS7njyFrbB6tyHfCsWNvVNbRw928+a
P0zx5k+s1XTn+kN7Ab/EtW4C8ZKIEIW/mLORhwWl8q4BDa7gbTlZzVtmE0D+82Rh
AiF8Vzz5HLFgTmxDL+hqtHoIOZNxfrG1keFqIaRkr+x5rbP8CUSUjxWSubngx7YZ
84O+5VH6kxSnTa11b9oMvEUNSWFS983vaXoBKjAy7zKSPWlsCvy4K9K/T1CYja4M
MQyEJYNwPWtkASRtU/2p9UFCd216I0qYxhBFennvygfPTiRnz5tS2brsLHnzA/zY
cdUR1hHgRcP8wSpQTJ/RKEjWJHXItQGIR1qLZZOvUjlF4BR96c90QYpSAHxr8Gqh
g6FdymjVUqYn2IobBR1QeTMJB6OkkH2J54YfJ7w1ckX9UL98eOEFRH+0qr3T4c/1
ZS0Ia/liQbEilZNnq8U8D3RM2Qz77N+eKNliABXMEbnymkmlPHVjwWL2WpeO8kvq
sK2DCOrGOVm4Sa+UX5fhCbtLHdp/jkDQH3HkIfSiueBZGhHvOeV/ygaGclutqBGL
WjZGRTTVKdDc0NMwdugObiNPXczJGwgMV0h0aCil/qrwzbEt9hUGAkYZcEVSPF80
wgXJF+xOXTa0UkDxtAsyBDXRhCnf6QMAp8SMg3kouhfFNr83SWPbNK6OC42vgfg3
cixQ/g3hTQ6ufY5kVvMgmC20Zn4r4TvoYJTS8a9Fr31p/8uGiQ8VtdPe5bAVhIOH
iRkn4rc6jFVeYy7Te/yk6I0Xs1DZGqjRsoWhshtTA7d3bCCNh5VVwOe23NadEecS
ZGK86oNKkLvs9obwVk6HUvrsDLGTJgBLojLqzWysJbhzdhYK3Ww5XuxIU3x2ZIQV
y7rf36RfXIhrOj81KZKMmCh5AVz7X4oNpN0gXGL/NNlJlUX8gjkTPMYlISFOVD6w
2VabHgfvH0gHL+Zrspxge3SwBMpvBdMZ4uNpIbogeWj6HcRajk3BAy3rNvKF8+Ui
qRoMnbpzPFgOrsteFui2vABsSl29P1nJq+aghCehDL8n33y/KeYfjVqJjZXCVGPH
/003E6K5xRqawEdqPmjUneuqgWEkzWbb0sH6INHl8+t/MsSGAB6jBGIAvG0Bwl8z
GNsZ/bji6SPFvYfyZLdviiMV8BSuzB2evO4gu9bzRNWvVUuz99sWJSep1XRt7UL4
BHogoElKba0JOK8nLO6Eo5ZKUFC7CQgx95S8Jq3EXDL2yzOU5BWB02i7Malf+L9c
nPhJow4N1GtGTsPanYnJ5hMsL7lsrXuKJev5yUHfYza+roN7wnlbXxDPNOZXFVhs
87pTSuJk6VDTn3Pappj9Z/FBVsjoO9xqtOogdyUFU0mTsaaDUFcraOGyrnY6s3s6
EBTtL4loXyDIq5DlKUdVNnH8rIqbB8wMLVwLQo62EkyyP4Ii6NL3VZA0LZ6hhP79
qSer5OI87DhUHGBx5RyuUKNv8I75liVoqxsoPbvFYRJxWTZhgp3Q/O3FDIRl4G+b
qiCCRP3edSwg5HjuxyYMn9oIyvwMqf1I1/rAgHsqEl6jVw9Ke2pA1ZqKLH4FAq6F
ETus0k8bpMUWs0gkSzWLAujaSq4LZ+NIMv8ktlQeSP6V5pdNNb9wI/dVHBrZz6mO
k5Y0Bsdp3//NAiSgqfaqAWNIO4aaUI4hx1EpT3wGcnm0p1uc9B7fVXmOD6JmL5D9
jAPsxwQB7JS9I4xmW9miEgcWM2OttdofitWhwjlR7/H/n1oTzag7b5m46g2g1GYz
gfTX/FC8JqpuVZf1hmCIYB8zTAlVHlpyV+/RncbYboPGKVaS9Ji8mjnbCdzoGB0m
5aZhoXHfplxr8osR+tJY6ErtNTOSHU8Tm33gIJI+qc70ikXdWhfrbqfKRLc9PwNn
t4643S1Z9clAIIwABQQX+BJT5cbwtsqNs1j+Oqz2AyKxgK5EU97Z2UYl8z8kcPp/
BJSpJCxzD3db6OnIa/dtefleoVBtYVMsJmaz1rcn02siSBiSFf+SrK9LTCZzUfOl
CGDNFNeIfxdAKDF8cEOLIpyoWdmGmnZQ2XG4V3JyLrLF/Ym+3eTWaURldnPjjvU1
HSUWETIsSZAJObDV4kHosaQ+i/OyzGSrORQpoRrIO7LbbDMYAMFuaLwgDNAUW7jV
1/bcqrAzVpZyTkW4+pHbDeUlrl8fgyJPN2xT0kZc+RmVrLYVz/zmJ2c15w9D97ar
s7VlniaQxsmaZ4Q4YVZq3m13d4NHeOWYBrp0soJsgO44VY7pmmk/a3CASpb2rb38
HUughn+uMdev2g5QG641j3XtQ4ak4DLyZfrJGdXOANuR8m+0DblfaOETGqa15VxN
5ZPdrBTr6MISPlEo4hXIXx6sY6dqehZwRY7G18lxGZPq2QJgBYxguZikd3fA7K5q
IDH5aWui+avu70BIyGBeqoTdqAIJk8zVyiErvW5Siri3ARUCEKcCfyNr1J3m5sme
G1QPYmsYVG77e2BZA9poDJ4+QCi5HV8mFhpS8lawpgw2bWX7PELpSh0WsZRBmYDw
ji8bXoEmwZ4sWrpWCaD/oFa4kgcfWNYXAAPrEOy5vqrfvjyJE1E15GSYrQ2yROVa
0EXtziiwEPkH89TJBSH2UL4EUNtKR6a0+icTlxIiCOCO8GSJffBgXQk/GjXpNV2Z
Laxn+jS28Wg4xSl0VC2npeGwaQyXZUcHZe7wqQWWgVSHltMgwQbrZnFUzsTz2Li6
/DQlYs0pJmc5JetdXLSKIN3zUI0WGJrGTWLQByHVGLDrN2qB26YabMOy1DpKTHQi
xC0Ptl67+peFDy4Be6DCUZCEba8mQF8XsMQhMRWYLIH5oOW9hE0jQVDjD+BU68SB
bT4VlKc9zfux5fcObhIXUcAwCAdWPzU+5zjQ5b3TCQYpKKPnHS7Dhj3YEJ/dihEY
fKE+LQSfXjs9OPd2MDJd2YY8InoEfinlndKGD3y+/j0LZ606351ZiNGeoOO8cvgl
1D2KIP8Ww8A1t1/lUWrSpaYCIInBrGS+HSOw6axReJAZovHFDgkaWa/O/UaIYbIM
I76tF9S/iHKuNJgrEahCzHW/S2BGOTmAFm/S0iwtODcNHgZ/UUTDaNVivE5p2UvX
cX9zSHHVUY0enoI5Rr/tuIvFWnwUDOcZrxTgwgMu4Tc94eoK4ACa0iLdu38ISUTM
Os6DPse1Pei4uaea7o6EbKEfOMlT0B0sK7lKlJjqenNiBW00nSkLt7VK6H0cJMg1
x/iUv3reBVlxWb5gf+vzPnm0Uy7cwszl18CdXO4wjpTb5ADLEvFwWhAoRP1VNK1E
RhRTQPNk1HdVSEmPbzM2j0GEwCfFzI0pmh7/OkJSHF01Q6R5uKRUfhuyJiQpyt88
cLs4PwmOa+bp330qu6DsF5jQjw/ZJ/KdEdXd6TbRHskoCpFpbRJ1YzXr/7aS3gvm
HfNHKGQ0PALKcDjA2n9Y19qqF+ye2OtOS29g1vE2T4nNnrQOSw25EDETWM6lCsJ1
9EGUVRUpCVT1Y1tR+9heEw7wUMaI8QOtbCenjEWsQ1hLig+Dk/XIJOC3xLEJI55+
e7VB6P7t6OfU45GeuWKTf2upDQGffKRJ7AIQgWuzjA0tZT9SroVuBy96pmsEz25v
GQN6wGfwzbMdqAjV9tEcNXzia5Fip5fh+LbhF/h/1J7KU7LhE+tMQPjRZ1ThKhut
d6/KkLkExsJxaSfEyXd8XNT6i7Q+hObsnn+RpSh7M9URDhpmSCFch/2Ycirs2GhS
sm3g6A4xvDnAAsibbHrrKUc752h8gty9EvV5X9cJoJZZMfiAyHC61ujLvaQXqltE
nmUpyu8LvxzwOsfacLjbgCUQYJ6v4d2HpFBE4t6SnKk5zqavteRy9NTINT5PEdZs
6SQpsAyTS4zQSpR4b+xzBlJgXZFTc/sA+Sn3oCkTcnxEP46XjEEHR+nrXM9oLsjU
MVu0wpR7PlnZOKo03G68LP75G/UkSR3btiYnZosCelLdQwhpzt3wdrVHc1Ao+NQR
o3NUe4+xF2Hmy6/vAl2tjXzEVmjIjWBxy+bkFKbtBCNaXdsS65qv+R3FTrfeHRq2
vEGQQtCZ98heSVA3ro+Rz+xwDZSg2mHIjH/sXebaigTXMP8etCaTIRuWtUd0p7Rm
WuipCzrhUE89Kqz158m7U5EeB/Ug7NDNj0d5ltU/1AJd6UWUjwWvDWXct40W4OtY
a6Y6KAhPOwWMxB/U/IXPctnl08Otk+u9XjQmPbFTFyhoEhztO6rTUDs3x+a5xWoj
9/Df/u5EZifpBUlB1jslsK+8H26tehbOah8/LU//BLjxlalfalVacxN5tGTqMuD1
u5qfCC7KCza71wqdCMGAl7Ng/Vty/wgdQ0xLUUQQ2BJwtcEfKf3u3BfAuJ0NSCqu
F1wdR2aLW4O/Zfhsr2MplpHAHOrzAQtL4exDCuMHgTU/r7fOQZnHFJoU7saWmTam
wl/h0I7E1p/ukVkiLWBl74tHSmHrwsjI0ysxsQVrfgMyePFiCio8IipHcLN/Xck6
LQ6zPVc91IxMsFeW0GjFv801obcO9VmwSOVpHIZP6sNZryR8MxyMFtlCqsc1jhrH
5LXJU30FoU+GJJcdAh3/i3rp5PTsy8ezx1kS/lCwlf5BBtgAcEJYZOBSdWB48Saa
mGtzLB8PPM7vdWRpnSUgGNtmNVUbpOwUIUmuH0BW9NDz+NlRa9ZwySyC8I7v/iFE
LMexDzQjW/5a00se6CDLofoterTIKefn3Esgg6bRonhaelPnt83+d0CjihdLTW7Z
g8N0DsdvoI0sZ5FehbriT7aNRbwV2vT3Ca7q2uQ+HWaKSdVP8hd4F5r5ncaQnkcn
r7dbCxVEB48ywnEQNrj0O2M/X/3zhmAP9rX1PAb3YlDr4rWRlReVsGeLDWnGI0s1
Pxh2TkvGqcw7u7+3KGyy9vzjVanrPgbWAMZ0osTelQeMvFFT5obELj0cX2KxeTLQ
+pGdKsz3YWfk7Ibnl/HaI9P2Z4WoS4ekJW711iFu++BndqAdV/O6sZ9JN4zvFpJt
X/3NGgc52lEn/5E6dcFPcT7Iq3n0AjF9n50lx6u5Z5AJN/G+puoLkWbQjO6/8e7E
tezGGArCo19wAMaj6DQnSrHAX20Uo1zi0/pMHVWe2cqpht285p4vZGcxEt+poxwc
eISFK0+l4nk7Q54VQzRyZJ4ACZVswC4y0IoRR6kU+sEaezUMsD7qEWkyMlonHon2
m6RidL0nHcp7h588d+hmlrgS5VAokE1oIcd0TryX3XnBUBqK4LQ7Nh+SoKK0L7vp
Vmbm6qT2hlqgZa6XJeqFMpAExtYHePD2LiznKoSf15ErQpzo7DYrP07YSaN6ktn8
PpgQGh1iGsK/RAUu20PiShJ8P3yPWvK0rDDwnXoe1Y37cFK+ZihcLEu8con+b5tZ
M04xDKBKf8YeZatyLQrR4hbyWCDvWqph7EuQEBwGhb+M/q/AYOc9s7ObDARmFQ0E
jLZ+a2pHYa1B4spZEAJPw8E83/S42Su/uVm6BdfEcvJYDWa00z3sfnVRHTGqSsUO
YHGByYndHK4wDPrO+mBg5wiBCyJLl1RFh2kQvUZvKpiwaoRkg5rUvk5nHDkN4FkL
pRwCMUwAJjca/pmL6sORySOyg/KKKzxSU+Xhl3RyHlSLKKd7vApZtIexxskxU5Cq
7W8ZcYmw+HP50KKyo2AuMYzWTfAMZLLUu/xy7gQ0uCOG2MlM2JilhgyNwKSKBjNL
wQR68B14dYd/fOSAj8sdtCOzytPnoCddV9kgHGoCabmu4K6uDwtPEZir7jqY5zuF
RbEUVmLaBjVdLlXGAKRtnEsGSIal4nE8XXMZhA66V3Hc/ZqIDHpPEmT42Bza0h3l
PetFtIN1Jf9QxmkbJnoloh8y8p1bg1y5fJ8r+JsyBe9m671Sev/L93wh/ELyXC98
HQfBXRAfu24OCkYNsDbioK98eNn23l/8PgK/kySyCAQUYWmyM5dnK5gKu0jKOWM8
ZdBs/hNv8RQj7dKVNVJK6OT19sALMdDI7DftquMAAcwdbfLbt3AgQfrZDTvzQ++c
SS4dTE1FWv6cPoLZ9ZtOGtkKth6eCZFjlLAaE57gAlGI1FJFGcfxtMvOwmmP+Fep
/s5wxUdHhJl6sVA9eQK8miuvCtxBSq/uCaw1ARzwF4JjfBdHs4TAedAEOTt6ax6n
IsTTQ44GwQp8mr7qrlyvDh5KS5tuWPbZLnTdlIzMK8g8mXptB/IZtI5GnHvngHSG
BdQfeL4N+cQVjRll2KFUkmlD/zSCVn0lomu5oCebWrJwXshVjtuhaHoMVJDyVccR
gnct99wTaRYKAl7aUvqj3M19/7wXV2fVQ9olnjmzNek/CzFt95TX3OYjwlze12Iw
x4JlNaxmeN9NsjwJUkGQaCe8t/R+is0Ur5s3iR39vzjBTN4sZtM5FZ7iuQhXEhYb
7M+Fxfi0ljLFHcJjLIGyBns4uay7xw1h366DdtE0vVtIWYHlfV9sN+q51Cmv+/6s
DBj0+0lY/4ZuwOSPFBFQmLNaJXjKhxXAwqqieqCIbv6PWCj+7rFjUr0+UXYdCp4i
93roxB1WC6wPB8Zf1SQ2R3nQc7+vn04uN8a2n8VFRoitHi2+6+5nueb1Fqj5p3/2
Z7z+xOQgDzuJO7eSyN7hJNZAAJV6duj8q+p3MT3faKw21afpEeBpJG7/Rf3F79LI
tHDiQYbc1TMF6yc6zG2TIRamVrvE5Vs5Pc5w77CDC8e9VKkjzpDzSvHRF56Q60FQ
7gt2UTuKoMhW/J9UGOypJ4oGetnGtgEn47JqEGV/SzjyD3V5yQhiZNzK5wvSQ9Uo
XGFntW8E2L+QEC1PkNtgNdMC9VuJAwKMEM89FQM/WKG4oDdKCAe8a0xEcnrAvqMd
Bm8ziBK+yS4ne8XZ6/jTCmxkJVkvGrlXNTF7X89V9A9DeAlllzk15ntIM2j6YzuA
PPw+xlzQPzYNFhjQ25zHaQRcSJWrxZC3N12LJrdKr9d4xld3pHOaQHC9gAyHnDWt
79zWEm8UagGZB+5/CzJI1Ah+Akd+001AKuoy/cJWL8mFRQ4xiuwmEzOWSqK4Zn3q
0Rkkg2m8G3ZWdiB/el/4JBOCnz3VS7mz6H++nY+FHXgQ8E5Qgho4GTLzO3GSN5iV
hmjDo92ou5z5qmDeSvSEjJFByDaDTVmJYPXVj8gOWVrqY3AeDqqrLo5EJhvTFGaS
WjLFx3DZXFdyK4/1SNoe3VYYnxkUxrnnsHaoQG1Olac779yP+9dzX4S/jedBkv1t
EZp8bezb3pvWUcf/6maftfufzKKnBiH10Mj6P7wrliegJYr0+xfAU0zhttuc1kqS
YUaMsDCEMwZ2i8Pq4Vc19Y1egDbuk5xhd/hosq1ndcWhh+9LwOk06nfonCtoNP3X
9ogMTsUGe7PReWUC3yLAi4SpRe+bCCnqksi3WFtT1VGwaARpnk8fYNC87MtobBWX
8x96FrITMvB7HmP9Toi8mL7fWfvKb+1r74c3z4IWdp0sk3wm6/lv+60XOzdgHjUh
1bWKHZjQJOE/RNQFeFfsU3BQm37JZenNPRCHDrz4auRzrlgL0KRq2jlPK+cAEZrY
PJnMYAzlKCVRhVG96s9pkv8vK7FHMCoJQpxljxk00Fo9Zaif5IFxVJA8/cn8E539
eAIyf/ZyK85xL/hn1f6SiwWwVew9apakcH7HWyWq2nYhw24SsRZur1+2kPdF6NF1
IjFXdoBL/in+V8tRx5J8bRlgJCK0L0V/CXhZRxkcVqXuRHLy4QG14/gzs9PPu/AS
t08y+S3iWkapMjdX4pxgqUucwh58/x7Hz3lcw90CP34GI3OtvnQXpQpIobxK6CWm
bCGPTSDxpfBTtn0nGp7ShmjNj71UCqAPWrVgAl04zmXbLcZ+cZ30Dh/BUqZztN0O
e4zSW1FOBVZLFesrkFJF9bppKxKfP+LqezadIfFhMZy+LvFpc7xX1AGEpqGS5lNi
uc0WaykP61Q3WX0qhWTQOsL7sCN3a+QXCiO/hlJD59Q3oHElM58BWn/nqamXn6CA
ttSINdsuBzH4EGktCQ974ZdXliBcYv3yVIHUvJU0kIJffOs3qvJrD7NCJtkVkvYf
rkbyOL7hEcSQYuouYEcDhEJ2xPzvRxymszYkocO1Y5XVapoB3jr05ooInA4UsXbX
rT4dFtlX4fakKkLN+u2BJ0qCCONeBGa++Ce7dlNxBQB1stQ13rVoJyyYLGP5ZeK1
FBffES1vsvimDJ+O52WW/GyQgCIcomQAEDpuS63GB0wsXM0XsaaeceunqGZl+/lQ
wpANC/nQO2y8AoJF/XlvBJmwMS1+h0/ygs/2l7tqzJ2HZJaG0YJPd7wU3w63ccLV
zkkSzkGHlPnQlzmZRg3P/zU7RVbNgBLVSV9O9Pcf1L0RDM85QndwgWpIfGh502hM
mtoywSH5OSnAZeY8dT1tZdBreAyTJBWoaBH0IdyeavPbp+LAc3z9e6d6ECEJBMzj
PoObflJF64t3uwuA3ClgbpT/OKblrp/5gAuA0AvH+cQ8nPODPSJLpT9FIe+6v4Ix
emJW+hqbTbxYE8zuTZwhQ6xmvWOKAsZLyzgzENO2x2Jl5v/HkRRRxaFoJ2xnq++k
qPSFnS1artkUnwNqt8rCgcPh/DZQZgbSWvN1ZingO0Bdf5Q8x4IHd1JZp75zCfND
vHOvvDA+SFf4oev5Js96gXnVdi+ESwFg2vNogiodW2CfOTocVoZpV8Zv0/sCbdDe
NwoMTXPOzQTOFVqLFhWr+Q3GgEpZGuuUigHSq5aL9uUvSS489tQC8fh3Apa6n6M4
TnP3TrJvB/Za+nXcfvF284IYQfVt3hF7eSsunUyKDqsei3KSWFtmVAEsUFQYZ06E
V/3AJJ6nHsNKT6P/PrPV8W5xaGAjohgph1J8/22uoo9mlMgFYwr+SRjiES44NwJm
fZ6X9lrURaVCC7N7FstGKCsUsOiBh3uZ5bt1DnHyC8x79Y3EX8ex1f82tU0B41qd
DE5uqSdfr8tTULiXAogBERN159okjijjdJv4fdtPlLi6p8vPHrb/6N0EANdsAzeA
nH+9ySDjvvUgs1wEbjbEQ+HRmA3WZonCPVMk8PRkvCVHaKux4e+/y7dpO8dEY/wG
X8ovztREZreTf2gb44TyCeF1Dvv1fyOY6MBNofxYwa4VsEMCzjfTIbDBa/JBJk2B
2RuKfbf9kqhsbWIuMZwtGCMZ99sWlqk2H/IlhV7dAmrwLpAdOPJgazmkJA6hLfIw
qL9ek6jhUPfUPP0nBMpAQE5A3KiogjvXBJBAevw7DyucOlRtb2VpaEISN6JbMZwO
/rSeRobe41q6SQ7bVmfNG4AUMTQVgsQRKkHObxc9R0HqXEy68pvLhLVoa4QUFOnf
gI4CV8svEwQWd20KlWspZ9WRl4tfuGrZ334rkjMI/ya/Dzn1n/7EgICNKiQMLk7+
o87YR35BImHfvzOFNIaPQZeKUx+tvFTB73gLjksUZVbt21JJF+J2VpCr+MWznieE
6tATQMbA6OmdlyTFCrAkT3yFwd6w8lMLf4cU7oNzuSn7ZA+kL6gyyO9FquZwUR4A
EPK4aLTmQ/RwkZwR2D1WcYmNqjn/FL+dph55KidRigzysO6vGgOaGptJYez2WolI
PpRjc84ZirVFiMsLpp5J4P45NLditKWNgnFHfyPjWlP8ULIvcsBt+pxxvXqUrrII
cceyMzVuF+2dTqRvjReWUhpx7yxbR21Op332bGJE/Pe5F0RxQDayyOSK/GdChO5m
+df7CEGtW1PrEYQzZGGwYR39scecADm6dcFst4eGIFMZnt2gGjIudheSXZO67iOQ
OYm9yhtVgwo5yhmlDa2aIheKNeccf8TGFwNd8YkXr1ILKTeljfhqyJhHE4RNY9Z8
f93X/sYh/pelKxmpXVmK7h68p01YBTZZDhyC18AboqAR1NiKfnXlBYVqsXhOOROj
hA8vZ4JDHiXc5GSnoq7qtbN/8m5FJb1wKQqIDDbyEw2BdPDOf4sKG1hg2cIdWmvf
bxkbpgD4Wo1o2NsCMXmo2Wb6A/uI2/uTH8woqAmj1qouUF+rk8CL3rczTvGBCttg
0oky1NKT6+a7Ct05jwLVWqp3r4AxfRGDtPDUbvwBzrvCY+JxEl798cdexFwI9T/4
mVt1MOVj4c3yMZu3lAwizvFwuWIfOZewyuVo4jvwWVaSb2Tvz4vlMnFokyCIU8ZX
3Uv5cTLd6XvbrKbIHPJaWOLgKXa4q01Bz3IlSPZLVIUS2wk2FAmtfkuCaoDAze+G
bEBIP1a2cX7+KO7+xaCl8CKe1N8tXcujBNH+2IZwinyQyUHCCZEKsmmwhoGMRxvD
oQ6LDR95l7uSENNcOgwiAO2VVSwynIdZ4vsjQMP6+TM+nREMdCsZgRbAGY6mohGb
Z6gjZO/VPoAv1Yajices+sxWJ8eC2nFDwzV9d52qIq5vBynU7fThjvNPlqGRPNBf
HVzIwCeH0Nc2nrVr5Bc+E6fxhV6zhkcJ4Z+YERmaFq2IXRQbF2rRSSYGVgmzjSzH
CupvIEYEtVx/UYPicr4PQaFi3qaTAK6tnBlVGhvpoC5mrL756g+1XZt9rS2HzIUa
5wbRKbw40PXpxVpINOjrVC6bHbaGswPBttq6XkG7ThkljR9SO5sY/U+7dkJZd4XZ
i/xJkvenXGnwzjRtWV8MKomFnjN9/sPWbPv07vci1ZQffrADmscMq1gxoqw+374x
uoBt2iyCTSv22Z00gdzs+4fbVufGZYETSKovrAh1iZo+ObHmSIREaNqvRIc3whDp
kNF05tCBfDdRoJc5ymJ/n+Z4/Juzo4ncvi/1ZF1O9Ayqaw+C0vrch4gDEXLxFuoi
w0qF3+DwfyA/oSu757hngnHwdLd08uhkndQu0Zas/z4UbgUwYqslnSWOOVzHJvWB
gNBUMNJAowp2j5d+dceLtCorjBTy6pTZ/cDTtIQtICrXsL7dI2IyGqt3Q9wSmac7
IzbL3JHPiKBG+wm6k/a6M0i2hNRikApq+r74iUox1vsp7OQQ3aWrK8s70oapTOBj
PkSq0rmrmHwGIv1V/ha+q6TNGgbACPicSyiMT7NbOKfpEGCwYqUNQbEA62noPF7T
cnp0KIEthwQsfrTwKQRTTg+YCRLt2r/Te2DWMmXkbN4Ze8b0ZCeYPxzEs6kFhCHt
FdBAEPfjV+l0U4aixnL6yOraMd+/xY1nkC1ywNYxgFRy9DcNj7ODgKzA29Gc+Px9
qcsjyXoDJLSp63ppCzzbb01i4RLoDEGu0OOAZYAhaZg90zRVa0CqEUtKfLqPCFB6
Y1C8bG5gZsnlTgwgtsrCT3Hha1UkGQaMD/ls56LvhhQwSDazJxxY/Ogar1lHcXTi
adqBvAAqqmYKReKR/cn3tMROJEH53qNhKQQCZw//YJweihPafZfPNu9My4W5siKG
KIiSSG74xo7x9/9eu3++BFLToFuEA0HI1J22TLnN4iHvn04wnH6/t71UqctaHugn
lDhEq1sh+/74KFiw2yAYXdGOCPNb7HZSyVb4QqaLWxNASVplz0IiuafFxg8/RRHQ
PbmycoUFNE4sJWs3JO4upKNhJTmrzBOj7hoYvlUdWlYIihboNMbXcEdp5sE0TYHv
+lQMAz/hfujXdq6ef1dwiX9EmF1s96N9iNpFtnoJX4zLRk2BPyied9zd9KEBlDx9
MIEJryY60whpb4HbpR/XHwAUzQwOaqMl/m0dp6mqXKVPgijoDBUa0xR/2U3TMF94
K05qSP21VFDMji+kqGtnNUTv7Okw6g4C6sEmYGESLB/O4FeyAnxffmG4l0M9daL0
4mtjWo8rkQSiyRBmxmP+nNnUkmrz+qgaPi1NdiNKHK7qmZPUFwlaezPtyDnHYBnw
cez0oCKjIG/woRel27Kt44wAWRpBigVBBGi0f5girU1KB0h4tGfTr25aBjZmGiVk
6jQ7I/Thh8gOdMk4ytWy8pR5Vg1PDVXTYQjOXeUr25e+XL6PeKRKrBut25xTWXm/
Bk+29YZ37HNNgVGstqs7PuUOaos2cYJcx5lHPX625tl3OexqBukcOuIuEIP1NDxt
HdbW8KWgfqtLD8o/EyZRJ2PxBiETnr2+1ThkVIdLF3yjqW3YwMOy3HD3xx6H5c0+
Z7WgXnys2rbBCEg9RNBxr8AnZmbAWM3xhlAX7mMbpSz/JYFGKZiIg2sSfSIrMdkX
jvEuayKY3l0YRUyl4Rfx74bEYuMNsBJkaJ8AN9NNSnddx+RENutWmM6Kz5Esk8Bi
Oh2/Wnnv2GolUhcfDt+rEim1eX0V9Ug5k9ny6gYbFEhpT+vIzQDUs7gmbB+jesLi
43m+qgiwVYM4UXKZlzXdgDQzHcFbiCIM7LRmaYWJkhLErtFEztIm4CMjCn2oA8Sq
yS1XJhmFANezxsRFr1zU6/tUGSwjQiPfagOiNdfbanOrWVSavaqR7uWjeLkedfpp
Q1WDK5MzTyOk555Kcn0Qv2Wj/PaDigGYLnMJgicVFsfjxos8C+r0BNkhVZUecVza
n0QuxFv/a3L2ZCW1OwtlDZl1fJA2z8DFCgrWGae3KL+2Gg81JEtqwlkn+b224lpa
4BarjonjuJSOHOo5hjWDf2oms8AP6BugBgKjf5zIsc+ydYXcp3iByPJXEXcVVit9
16FgpfDTEp++zBQCUA/dBAA2qkUVtLYGryc7Vqli9plRMp3pexJhjQkcNxryhAPi
bArtq+GimVlpBDwq5N7E/7AnkBm4fMRKBkxiOphi2dtsz5RFwYYCL+Lqz2raTBHz
Xc+kGLoSkgHH7y5shgEKQO/OyUF3yveYtfpKK3V9dkNXLnfQ6HQ6f9R/drcNIXHK
Rr7SO8+aeWyNhvf9JaWjZRn2arOF4j9Z2jKZkm5fgzazC7RTn9/Ft1u0l29Es3GK
HEXF+kEjajib4/oRK69ko7gEChuyhFOTK/OgkXkgt6HtQrUPtQroqxxL98BhhxIZ
wD36rgR3QQxxNuVK2xOXN2+KGbWfP9Gy7uysxbJHzfYOr3+1vU8ji+IMuZzV0y6k
P/7rJbsRnMra6PyK9zPJYIuF5PTM15Z3+J63o6+QN3ZE5690lVDJZT+JsXU50ysj
fLYQ3F5lxIJ9n+TIMm5Uod2tr2dTBNAnXJV9EnaQvMtVwxf3tkhNV4V8THZxslOB
xSfrGp991BOplUsnpPZPWEtOnMzU94kFa44swAoVyTFoG8DoElnsqNDQAfZoXP+Z
LxIhozfqAOcHzbhwK0/LFW+Hifxd+peOp0WQF45Tzxe91IZ1RAarhZbgjX1XzamB
Ne4+G1t/6nW5CQjve8QS2t8Ecdkq/WrbeU2Q2sutt2ZXZDic4PDsLnA1yvpH/L2i
LkKMDTO14OlJMp3o0p1LTbkhYEeyGRcaEELXrMt2ndwyDgdTXHrfOSpxgRsfT83Y
BqgeWz4JVfT6aXj7Q8d2CIgG/nyc8qg7tqYwAAYCbBHCa+YyPpJmVamwhn0qF6E2
KeNUaxjLMO19vOLSmdZ1RJFGT1LGPuuEzmvX/K8WGRrLKD3ihnTjxXxbs2xYGrXu
K7YiIcQSAC1kQy++JG7MjL/3ZJBd1dZa8CEm1fgI7NDsT/Lt0hXCkpeUOxUJGiOK
CiMJ7BMELJ8YcLr9H+ujtnWQEiBuChFRohjR/43ssabCz/b4b4gah5u/lmlilvYb
dLX4QkrAJe83/2cDOpJg21l1f3pPSv9L8maW47FfY7pUGF7nNEKYNcZ/J6xWkC8v
sfq38oY5KsoINLI4KnoIy6xIaHArLao/ufSRDHrsf12tKv2RE/FouDVGnNVnYS+2
SrlR9wZKsfWcSI4VlqPsjcKOjN56R47sFCjfCIdXQzyePvjhUAM9oQPElFimnE7h
yVpf/hbKlcTxnOriFY7SVrFgxVYY/4ucmkX737MtiHyFD4Bx7osn1S/Byou6Qc7S
cyrYSgFJ8vEVmKeIe6Al+Qn21PJhJ5zwJ0rN8df2C6weRJ4NLWhNMMaD/wtluV9E
TzH9UAXkY8Lw46dLy5Nfh2BR1dGpZJ6m1r6awX6BRaDiC0WGft6WYJHKw/doyM6v
dXcmFxT/SfU8Q7toCABNo0Jdp0cCajkrL3Hsdob6NfFYQQrapQ1Ch3wTPKgjyoPr
QjUwmjMb/sEdLvcgNdO8XQEFH42DFwNRRPc2Nf213/fHCf87WJKV2jsZl7qRaXcR
oH5mfO/DRoe+Tlo5QZz2N2/m/MF/5gNAb0pxtKz/1pU+LVzrglrqHEkLySWFVZd0
3UtUqIAQCy8AgFEKGT7axUFLzaKrk5B81dfr7o7/33YKobaf9hIIDdI9GmV8o5DI
ee891zBvKWX8w4pmFCuEg6nXHBG3AU1xSgLmf8s4VpQFGCoxIHPsire5kBeZOP/M
PkQQE7jKhY9SE3gDjiQJfcV3n0Um8XvYkHO9EesYdZOKQVjkU2wF5EhVCIwinccz
ILW6ZICasLboevZIiVHM9I9XPt1XUr+Vz0Vj6tC+BI67OsctWKZ1U8aSF0eo/yHC
a363VGKbA0b+KLb3NKTp6z/sJtSdIzTPdut74zZj3ig5Jvbr6dPCU29xKwegiQCm
T3WSE0Xch3ybL3BcMxoqfMNZjvpu7z30+4VdD/7p/7yQxTMYxKJQakAmRrTmC2oF
dlFd21YGQVYZnRcRf+Og7ZbBB9jS9dkAvj3aA2fV2g2/3T9QaMZXs5XoNmCaNxWv
G5l/ZlW6zYC2yV68GE5MHrS9YLq+PQAHydo6vUhBosuitIzdGE0CnH1sypqHpW5p
6zA0oX/TvfOGtZ077Qm2Ex50Xkb9I371mmFqdLQT0rzOFuWYgDtPuTcZNjxQfysy
0x/XoP5FnGbXu9+/Z1LqW+RnzEqLRjYr2vIspOz0X3QYVzMS5EjXqOsKgvE29Jy5
VOOsi6YkIuV8Dx2Wt5qlEKUfh5e9AZJucG+kWTuNGq1KsyrZU1LfEPd/wiuE2oHs
ybdPqqduJKhckdFHlhIYIfiykBcIbge8GH9P71+N3BNgZM7qyS/Mm3YgvQ3yZqD/
DzEoPnuxVGCizD/1LsO2Q7T+BuSKybuSWdYB/yoJ3w9x/Y8RTgxqQpcBu9m1Tk9O
yxnY7Pf6gjCeeE037ORSeqL7DphlN9Pwfibm7xTlUAFYOWiBLU1IfBh46mH39+AV
be4NHWuqWZylEBkc+Fkg1VxT09FdAocPRpCCyF4yXDLhrc36HJ22wtVASwxx/6Ma
JYVCOovHCPV73HdV+IYkMgsLaYOSEpUh7NwiylZAJZWCkCg8YHA3LCj7bLMmc3Nd
TrSohSoSadzXr8mGkV57/QDdfRlTwvYjeSXd+wQb/TbeJwOYNp6og5JnVpCkDsF9
38QAMfGPiHnv+2Jpj4byFTgARQid4cROdnnKod8A3MsaPWi2qy5gRlQjvgd8FHMl
g79elrg9/wbCQHVLlwj4VWbO8aL6GQCyk86yM12y9Olag4d5ymNhMMWhoQx9Fr5t
HBgYOK3DDXmX6QC60Zn4/AacOiNVGjQDztzoJfToPNhyk5R7j+7agFsibxjTI/md
SXC6QArKTvm6tC9fnBG+vFbRC0boRYXKRf0Yi2tajIZYn6S+0D6I6oKjPDKqkni+
uSDwTXKx+MGFdxAisJb4HFE9Ywx9s7IZ01GmBihY3uM8DaUDJdVCNjswiOR3oIhM
r+XpYsCsXJZ2duwZbXombXOTRmSjB1nBVLeMGqZWsVrnicvtNzSUeBk2n5T0ILaB
wa7hVsKTY/mh90LgdaffuSOtTMpIbpdLlld03x13+cnuzSDUCLMUFo2NTEiW3WKo
O0QeJlwyP5OCp9RqCwY1TJR4ynSfKa66wcz5pudG9lKFYqd+MoA6WXtEcKYy7rcU
fkBzIpvyXVW1/gmuHIxV1O/ZKVtyLhWiKnz3tJ9tgaNl0yhEU5+cx3zsmxxs2M1L
eu9f01awu4J/O7e651640czRb0WJ4taRxCtLyxptzHn614osKdwjV13aNZrE/DAk
jXObRRT3oJ1Ue7N0p2LY2sagoJe9fvrQMzpYq0XbunnXw6Wb54TpPXTBoLR5/dEY
xZoBGM3+sC+n11gXcxUFotpEDyABKQfbYewOT2ElCFEJxBLAXJRxovvcAaF4bXrA
39JGu9Xu/UE/dF+KKicL7mm2Jx3FG28vKDgZ8C7qzORTPRNFnI94mPFAV1yvoVU4
96ggh5/8cZvAb5OL+PxINYTRq5UUrsBpdW4quCDjyQvDNQsJMZH9E44HkGj/MeJ7
i1OT0IQ80qWvMucx4HNIYvpj4bPgKSem4uXFGTKw/7hPGMrCQJkd5z8fMhgwmoqG
uz17fXOn/aNiXFWRhMEF/YXiQJ3sUYp5WXdVNxRkce9bPdbTSeeE7e0EfTUJqVD4
z/E8XU0d+eQOmbXuTE+6iNQleWQslvSiRc3lapJ66g/3dZENsStpQw1FNNEzBOc6
NfOGu1N7xoYXxLH8cqB5v4Mt5r6w5m/DQls8UPMW70YETy082InTU66WoeXO046Q
0zKOCZXbRUX3mj/ECejBgNsbJvzz7MpCQF7SyWYQnj50uUE6VtRmXbhewjJy+OnS
W21v43bh/gxCK6HF7FWD3fEBD6zGT7m09i6VAYUzYxw7QiSOB11vnjCWnuiTmpyU
TaPBsUwNx08S5UJdslWhKwnM0TQkfSs/s8PMEXBY7crHr1u7k6M6SEUDVG3hpmSv
IXG8JNnHZdTxZCElEf5rnhI0S2W6HseUgHfCV6USHKiOuM5XORuCQvzPvAVZXjTQ
Eiwoy0vIfluFDiBPzMT1kOu4MHSo6ewg8KJPIps8lbcpMZRqYmhFU3D3Z9Ey7ORv
mtW0/lmPQgaCntZlBK8U8GZ9rIAR40+QiaVblBnoP7ljY8KRXAwo7HLv/r644VA6
9XON9fb4pghmL8pBwIWEJKBHOC4mlqedlIPsvJXnz+xQvRdrkZ+cQ4OLXmZtj+kL
TJcqw9WdN+qnLyzkpD8LrAce98ZnZMDv7IvdCmaTvvDcdTeoJ3yyElCVWsO4c4NA
2cip+5N7+AF9kEBegc7FTviu5BXi7Xtv6OkQ6iTMWueHJ2gGWkgPXd8YXyj+hLgt
OnSlDUimSxggj6u+QDNfVady9vLvb4BWaTwxkFmU0NCv0G7FVovDBpNlH91my8IN
Nn0MXGejht1i/Mmq8+ymc7/xLWOzHZzGNy22+uuXyLuFL91ZWui9AdQwqIVsLmie
WTTWR7TXOPidLO1PHXO7V69vsZK6zlpe7c2uzCx6X90kRQDB8m/qepXUEpW2PlGR
halkGL7QOQyYcIgkJ2LWW2YneJxFFz7OqreoRDWH5Obh+j3cVtqQekT/iopu//OA
gFKf2NUKUhyT3UztonwPTcOuLdjA5wg4U6Q4RFaJvzdi5nBWK4Zl9F+w4fJJ1Zlk
wSsbb2RisiybA5RZwqNLChNFrTZLTSYVCe5sE5zyoBQxoidF/dYsYVbUVuUZ7vMu
06FeaQsQyg/UhSGfX31td58u4HA01J6xSeclT6e5Y4dwCSqwKWMR7WxCeBxZYCV8
6oW6FGP5Xs2a6EdX3OvAkXZrNt8dJRhRJfCH/itj/N84YPs5tCheh+yvP4CGyWd3
BoDSpr33ylazZwmsenGhOrG0Jmr7X2qapH/HZMqzQH0CNnG77gNrmReFchTS7Qhp
6If7jYlhPRUMFJ6Ci7vZuIX03JiADrUWx7zQJDs57aLGs2kj9B77RsCUTHveFyPl
THqqBCk5Te7x058Hy1x4mwb4wwXFTwn53EYyf7uyZR63i9Lw1Ia6eC6e5BIuYsKs
dfL4rfsNc6jPuFAuMfZY6Y/hzPQc0pptoAs2QUJXnI+C1oezXnsNW5Tpe22CbtyF
Kgj9M571mEUEfUih6mvSDQitbJWfHwmNGzX+bnjVIqkVy3Pax+G6vUN3WZxDY1/j
eACjHOJndP3wiHDqsaytU+yJY0dCBMTHOR9p3qV3DHs6KWfDgIYPSDzKtiF3wY+Z
kka8PfulG4jtPmi5pupM18hvonENwiUppAbEsN5YT4Cs1DbT8YYbIqlEliFp91Ma
zSTzuTHAC+yMhz5Yld0PT9XiLb+JWn5jrbdGRaAbSINodIggLmzHasstRRAzRQgo
BKuwK/aLV8XZjA+CGwPxFBTrlCo/KQMCytlORmZv4AA3t16swaD6QbUh4Jbr0Qm0
7FdAztOaLkrohEcEeJWSkirVtDhh7IJh6AElxj/MHPmfe4YbtpZsxR81nn4vVrD6
3Wlyo//7IDi5Jh0/dsDYzuIR5xnoGzD8hPvVvIRjX+0Edv3gwH8TiA8m+Lge+ELM
6VqTpyRwEAHWYPgM5CMJF/X+L+VHYgdlb1Bn42WHCna4og773ydq3yUyQFP1yPUs
OEqjl2GS8CkfY8fetx7aLWDG0KNrPFTd9yC6+rQsmuIQiN3aZbxleAxsPuiOpswZ
6DoZybrkOQCdCxnMTzHp9yLYAOp3b9vH4dJ9+4RJvAmyzP5mLxJM2f/9WOJsfn3i
Pv2rjwTDn4MdYEVj/I7HhCERzQ2n1BpXBm6pP8ufmXmFZxJjA7DnSIwc/TMN5bcm
NxX75ZB5rYNpwlqDR086J1tbxf0UbgH+hZ5ZsXKi70ozDRSXr7VGBHpz1oWjtzkT
8hSqjsNfx7rXhQl6OrpoZkGhpsC7WJkv6QZCLlum+AIqFUA2OyTsY/yeZfi8yFk4
mRwOCTM+iFZFxh0I542HccGvUzCK5LfCiY13kKLD6VDTpZgpzy2+lIVGK95qha1x
26X1xzELB0X8OFCD1FMqzhzm7UQQ+Ehps1EWo5O3rzresdwbsMKSsliF4Xudbw+2
bQVaKvanRIdXhS1UnZEHu3f6zrXo9h0l73QQawxZDJTNMXo7ayquuGzuXKlJI9LO
WydhCGDf5G3IUAefEvHyXKtFFQ6LHO5+d8TtEcyGJT6qlt6OY6w7P4xPYQ+1q4be
ZlndYcyNnphNKLDJDhMNXu1Q5LVolfDwVIAXPxVCanTy2UFy86Y3Ha74kxxpM2gh
29RGhAvQkbq0U+O9xlpbFkafK4ZDqmBHszQsSJ/jBADlCkXC1uTu0gWnnG4lJsdv
iEWIkUxNSUaijeYtGIDTwDS/NcKcuYMuNpwZwp2EVeDgtFqGyTkTo09n3ef3QpBN
2dP388MAt3Kv6YBSvK9rI/XZkBdm6crkL5MoHI/xvRQwwRh5bl4Q2cyM1qCUKXxA
ERn1rRoq/iXd/ZBg527a7djM1Mls08VT87RzOuGPsXAwod7GJNuCSPN2MYIlvFAH
xSVH7YTtIUqDkGcaWmbdoOGSHuo3A5xFdWPN4/Z2cFYqQfNOlGLrvZLI9S5ViN44
puU9IdcnF0JkUJ5+3veFtruqpuaWd2As03kF/iINFxpJsGeirhbFdJHOV3QkbDsx
NQqqRFcDAD7E4RWU7T7c68l7cobmNCB7AK1ymVTlX3i8EZ6mQ+y5ha08JkGmJ3H2
YerrnBjt3nOd9npJqqCu0++KZZFHdeMLMD16Ko5e5PbgC/rWfcxQqSC4d/K9C7N3
x8zCRhAiDwZnnJ50OVLhX2dH9tBUYUSrjlkYPi25nal/tFE3lnuFBz/lsso/o9Nr
kQTx3B9kRuZ+Az9SQsdC29blzad5zfMn2I9hJuPIabG8NlDJvHAn3Hm2aYfSn+hl
E2S6GfUjs416Pze2JFQ1FeUeroNDkrTr93xGz22iLak8yZWXXpxKNKpBaHoTecql
AIRFMy0XA9CkhKEhAamufnjPwgeWNhS5e7Jkg8qxFqeknBPvkgs4HzZ45JNiiCkL
fG2hLpiRbA8MlxA6ivJTwxxLthg0w3MM8wo3+kRlsfYDBG2UaW/0sM0AMKH/hz/q
yUSl57TSbgNpAk61j1fM1j5RX9664szbEIXgRoy5peqiZcwXY8v6uUz/2W8ROPL1
8m8kgGofeISGaE4I7QOoZ0ibHeGwlg/8isyfOSOISWaXiR7hNgT5mPa6Ig/VBuwO
FsDEkP5QyrSFM3KgigEk5QgxGyzmuN0seISS9QQJZrzAPG5zxmjnQMxczqFCjl5t
DWN+tLpvbD1BzteBVpNMRI68DUrh4tEtoQqh92LaOPT+EHFymWqhoD0uSzuG3hmA
X27d/WwjHrax9bAvaDwSxvMn+LGdIdcBl88zBnass1+YwE478w4KllzF+re8AAZt
Xzqi5cCuhEWO7XA11HMVqF1K/XhWLdkKbautdFLujZd5nRRkIUdNsuAxWVxCRhme
PQ8r/FFZmOJyNi7al3Ovn5Ulp85KEUs3rYtPsy4kdu1eoK+HU+WkR14voRYvrd+8
/Bnl1bkYefqi0q8R0sMuICpu22xAR6VO4KP6o0aFlOEyN/aNDSFy/vHoW+3aE/8d
ej6LNLxp7SnE76E7BCyzWnFgHOGmeTV0wqZ8qn7dEvQi5mH1ptjw2c4XikR0Sf5w
zE3N9wZoDJlwLPoEFXxboL6NioiKEGuG2D5TQnjhpzpwSeKeRJs2bvEv75uLS4Nj
PGFtZelz4sZYa/TZbBtLMAoRWdKvd3hPURhKmO0cbUFNp2ObQW3lbSNnjlkW+H6L
PESxmDanM7Q89dYsWOxWjrfTHO5UOoGbIFOQov54Y8m0qUGj5cTm0vSWWIM92vWl
JoDEcWDjODasI6Qb/3Tt2DpGYKgYWJcc/N/N8rRIfPjvmqKMwjHFmZ0T+JnaJEkG
aKchgu1A53S3hkAqg6nVZDziUk4Fr2c85fUq4k+hq0wadNWxZEH9wSLjNvcM5QZX
R28vaxCfBESv98WmjhTd2nb0itc+muhV5anDlNgyBxtTBIuaBwV8Qly6+3Y9G/xt
TkUN2UG7NXPFmjoR8tjxt+Viml6Um78QUJ5lP8gr4WTw8jrJMqN8VKZUAFZwsqYJ
Rc6Zl1VqQ9Fu/ISTXy7Gh/9QH/oQd4TY9wwWF4AiHwBoWnckgbM1JrP7Oa+UtP+E
KMZiQooXOL47kkA7uEKBNP8V0Ieen81Rdh3lk42W5gqe46L7dEYFEmfIseZQn4is
Uvu17inCkPMtnN4x/ZurRf1GD1ED1h/r7L9lcEXOjgwwx2lR6yEEsHVyHn5kaOEH
pbVQ8HaiOeNsCnyBDFejRjJjPwwaDzrGkxeidG0edkIhxhbiVFq7zVLbh+X3ID2d
UgwXhcLhhBIqtpBTiiRYy7D20oKlukfvLxsXPjoM14F3CBqG/G9se5ekMdw7rqcP
NzYfGG449MPktYflS/U3b+MY3Y+0vu3DlTcmlUBKH+uxvqyuclLNLGpRYdxXgtvb
mMWXUlJKUYf6o5S260bqvSlKaBCrbDqcY761xG2ks989jWqop7+GnZHqu8uhrr18
0VZmdTzMs6arntd+O2nA6rI7tWeorI5wEbrOFSnNe6uYwfRnQduhTWrHtrlxHWWx
KE4AJ1YncjhILpT0FW1hPYcqvwTq1bqljK8TYl22aiTC4odLYgxhRxDrbA8WqIhG
T7b9aEkfziZ1u+DAhv3oCSi7o+e9/1p9QM2iSR1DD1SZJNEybZRe9CENDQHt3j33
om0w8i73ieQi/KKBUf5Gq37XRIvMLex5XVMBHQ9zFAN4Yerr50jQd5BaDvil34XX
k1+qrHfknxydooy1HlB63pvIcQJN/dttUjA50Ze2+nVfzDEdVoRD8G0I7TCqql0W
mqhqcxI1ryL8zmxG4Ewh7wNKIM7MP/x5pn25pZk+hHAJiJozD4N7i4T8CQ/ee8gu
H1PE1YpzD/NahwjjUfTgkoBlro350a4CyC0x7tdrftxB2zW99ScmVKlpp6sFMlVd
Q2ItP6/dtGhlUuA2MiUczPmmA0giGJ5wSQeUhdjha1VWUW8yxvFi9TzOJpSog+rX
bKBP6lzgxGx8adyyizHSZ3PkMcdRXMDsVQgNDk0vzVNByT2RxUJCXfbgGdqTNXVS
BSSjV+WrAM6bI6JQxPdapLTPgi1VagLxgyUhyFVGpvdV1FZNUaqJzrnGPJIOPP7Z
ySfQEQEIlaqQCOj6Js86vmZcx26d6VLWokuwtR/rw055vueRuQ+iEJcMrYkqTSr5
LhiniNw0gjJaMFw9iKwUp27qwid7tjPhXDcCsk4s5ww/jy1UMCE0gQNzCcCVzYgS
v1ZlnYpzH6DIaP05HtCDrETLvjVL5qVycKhcx4KNIuJJkzRQGcrNcjZ0bwkljEEK
aLt+46z6XYzZmU7FgV6n4MeGVXkhGl2mLRoc1Yr0EtYQDcYHrvlERFe3jpar50gM
RXRX4pSiTgd1nzQ2mn7UqupUjxIv/AzoqF3VwDEGu7lQcbN2AwslXOcf2V0yJLCv
wTyJLa7lyQo1KDABSroBQHmadW/MhHqPl/ypFjH3D7os6QOA7x+z1jQsQxB/zZel
/j7Uqc8zpF+okxTg8HlL1duW6xXAz5WDe8mHiQqbNMKZ7xl/f1qQMWwb1hnJdOLh
EF/wBNh67I7YTxP16O7uT8tOgvULLQ/zSX0eOOQakCQGxPg+0L1+vd+9gK1SDOYk
fDb7EnBmA0NuHk1r0gMfNLbjdS+a5UD+b2efs4E6STQnJymPrkTehFCOgNY1IBjG
Q1J1V5yjQ0P7LrNLUxOYBKUjp3/3PngTnecGHNEGp8THimFt2obM/Mp/MEXuxRGe
V3cOEts1kg3xHGNUpQL1E9ulspE5DmGorIgHg2LcFuRGhvgaRz7Ho7ZYdKqISmmT
ppA8nLi37QoNdwqA8iKhF97khzBD//xov+JnlvctwQ5AQcbEQLGJRuQPx6sntLDC
LwpzVxGP92vFjw04S663ZL6GUEnUqm03rDiDrFJqq9VgffOV0RF06uUnSnU78qrK
xYaY77b+tJEQtTUX09Z6Q84uhEWKvWZs6yLVx3aQh9fFsKxddWa7v8mH4K+R1Opq
MSiM0rU/9nehD0W06oTVJfRIheJD0ZuR7jOxz7d4ePEJcwcdE/GURKsmcG0IYFkc
VQUwSF+/J8ZHTNVZ8MKK45LaYvsVpO1V+lt+sl3GftEOzxXpX6BxVYJaes6qUdXK
QUOeWuUR9Ix3sC7U5wfgGybepMqltIf6nFkrZgzNdimHuoGbfSMFoXnkXJzXmOu0
rvmQHaxNppC2jI7IanaDiArLubQ5nStqW8Vm+S1Mw8BWoZiV5DpT7HuTO5DGR6cT
zcrj2LGFYSdgstEilo2eDTYx8G8JWchpdQrI1bmLyU0Cflzd/uGwCuyJTyHY6pSu
NbcV07fICk4pWb1700MhITrivV8uHDjkMGDcxlnPNgU2rgaU9TSV2fUoXNv3mcLo
dFpW5bMn7/iz4TYabHdnTQnkjA9Af/EhQfj9JFdrxxjcPnVgg8orCMLRJNpwFjQd
f8htx0kHbAtCsXFW0f6rmT7j2HF6s/NdBZSINI8fjYhEn4JYTZ1o5UU5UyeSq5MD
OY6nrR0bO5059gGLIqw5wPJLH42V2YgvknqRvTI5/8AdfAnROpXbU/cvvNrCiOr7
s+3njtWvnFl1GStQEFDaRDc8oKdWMhOF/abEnHqL4JSmnE6PFXEnWXPFpcR0aAXx
+QWPPBALZIVv+vXFiuzXftyUEjDBb5d6YAWXNWPN0RPHdfmXf8LgAYXtaUbHCL5t
UgJIFE9g+22WOcLdW/aIMgLQn4Qkjvpge3PggcQjj8U5NsZNOfyFbLGrWzwUgW7w
PLR5F760bLXNgwSHjnK06jJs59qDrw2wV6ySiucg4JJbrdiIYre0/ozMtDZNZait
VXRq2wITjIgVF3oH7lGTCuRsgnBzs76qDnSsdN7bQNHrQ80v7cqeyAlk3uL/QdTK
sJqz94liL+Jar/VCW1zmk/c08z/HM0SB15EPkTYHpb93Df0DRNRJy1FUszyxuKoi
7iLqttjd6Y6zNDAq2QXoEsBhbx+6X7WY1YguaNwpQ6z9pCOrhTK0IgRil3o+kgCw
6fYZ3J9X/PR7jsFdY2HCzloQntptFHTP1Qen++3Pl36RchVgmp4b6+1SaPNT7XQ3
ubhjLgUY10Tah1ZL3yAKcKRQpC081jIWSWujCvf/mIaZyNm7sHhFnBL5bXnqdsR6
mpa6NGbdfxwfEL9xYn+T7ZFdX6s2SS4tV9SR8X9HRwsX/0l6E0VdahEZAOfBun3l
hoIbiFyLO1tRhDqka8uudvrbrP4wxudSSRWehK2S2hEFGouSRhVA9/skZRzNRVgy
ReQCx10hmTSNS7o1wGhIhHdAncn2ibv2lPm0NJZ5IRcINiU9nz8S+2dHOPE5uTgB
nEeJdoFLSrp5l0sJ5qRcKeONOI/bYFnIUADFiWiiCDQf9+O7s/b+z48pPji4y+Se
SGtmdnEW3lgdX7jxDCsutZDmDxbz9P3RGDKjJMFz0AwdBvt9hdDEYtSm++xTB85O
h4KwVRT2Xe/AOTk16A5txrCbZSYgC35d42BI+g1JFekvhB/sV03a/PRXgalh20O2
/BAS0IAr2T/0PKLcfPFmEYLsZBsZ55yfM7+dVKE6zu5NKaCom4BdHmCP596baHjX
KIYeDK/x4PgPG6UfhDh+1DcmeV4rQFdGOB2G9Qu/DBWu/1ZpD2uqWGihXzz8ZVbK
ihZIuBMMq95IfgIdliR9IO80Du2/4m5JtW+AzkKdmMVNGWeQZ1KF+SepnGNX/XnQ
WOiiysul3j9DCbxsKV0EFlhI798WrU2WoNxxh7KeD8xKNLqAwE0EqXl66GwCsj/h
g29VVlRzGW6KkwC9otXmwsRAHrXB0fr/c1qaenDG7MWadPks89VWH3sfFH9eJHP8
/f8AMSzB+Ei4nj9ZKM3i21zv3OKCUrKmaOr6JczwWj49w2PgKC33TiGBSstwo+MG
6+dJPX/B1kE9miZi4eUSJz81DCX1PlwR3TEVlZ7HyTRux0RN495Q+o4p3l0Uv1N5
Fwysadi83yA7aAETws8v3rFiEjJ6RoVfo6K5FqWAeXh0MY7VihnwPGlfTiI0/7Ri
ZioeohjpgxZeEHbb6xzKGtwGHkqC7JkcQpPyGwUFuBxZupz+WqMUxGcp0cDExiZw
nJ44j625mUVifmFKqAS9cnCVtHyUt+/sNL44RNSVSz9CKqGeJvZv2e3o1lU50xiS
/bVhZC2B6BONbGzg3k8mJZFzOYksQTWG9eHFb8btD6UtdQqde/pHTrKHaguaRU0b
oUrHRPj635h6lRGSVHInsHBsa8yj1OBA2fsnyigXW22IjuHUunHFnisAs5paFPuQ
5RMYIx/IjtOjAPTlLMjLX1rC9QdzeaTF5wOyFwtClbLWzBqdgiRlBg7htQClwIzV
wTCxOzSwQTSGVdXrrAPn+/lxX0iCDtC0HIiOBTfArZu4t3DiRsaFkArhaV/4Khb0
AA2Ab2OrfilnEjyiOFSg/RauOEt23tXNUMU9n06qrDUN4ubv9n7Rw6EDIrE4AIm2
EDg+C4OfeODkoAv1K+25SHkEAaQiSL09WNU04Q6+XNcIfA/nWqui6Uh3Bbpd0YMj
4/InQ/VTyvb6HnD0RalvcZ4W6+8HX2vQzy8lPTtABzUPpHubG8aFlaEB/7hlVWqx
1Gu8UloNf6bMzKtDnN+AtPAxaw7sfTbcMBlyU0pphTDxKsuqgA5UBDxA24U+At6O
O2OaUh1f+sXjgtEUeRvPIrPC7kHqGSUeIw/Byzt2e2DRwbQYWPrRObEv/O0wGbLa
qu/EEL3uMx0xLrt6sUZUVbrc6HgdDYBYE23k597iMvYtpbxgy5NmhXsYmuROLWQa
iAwaAdXDuOhpPT/9aZbRw1qWgl5GaW4E5BAE/FRkLtIC7wp1TL4fHMCJWGJoubHp
WKww+dbM0iFc5tBhU9L2Ru9V173Zs7U/kXmqTHm5KB1lyP9p37YpY2MQBLSh42Sr
+ory/HwS5NZ4EaqrT/06FveY0Q/zS0rdmJbtvHLF5KlZUxYy3CouBG/s6dDdOHEo
V+1B3W4gPOvlecqHL/acux6qPWBj7+shWZP5NPNA91Smvg8+Bf2lxq/6IgSMct34
mDD5i4417ChFuHo8WLHIYhSQhQjp6nb81pnhKi6Wzv404lMPlV10wn6DKe9kPpKv
RK6trZ7XnS8peJv9oIvl70DOa0IKsQpjTfG6ggOpTjBffOs+rngpeaP1C544pv/i
OyjEfl6+NpdrmCuMrx/hRX7HvApY+Ksl84qKw03cSkuddgJW4p9thwRxggVu9hvv
GzpA69emQ4R/sHp/wdHLFmB9HLSCDy505c17+RBY9KLnkYTLoN1tayMM0CT5iPjM
GLcbftqt/EQQiiXqnE2rwKWZ5aoM/I7YeE2aUVhywSoj/7KVP+FIR39qjv2dtK6+
wWDFH4tOJDk6mtmQrgcK5oWf0+9zD0Ui6uJOyPKjaR0ZX3nxqYwc8NuD3Xci7Skh
BSqKX+WvFTBm1pr5ZMq62tlPaA/bCzBgGVAEEpbaA7aBo6Xa3x/x7uBXj2P+LxYp
El96roVcp/18TFjEQH48npEXFWOZ3UARUQ6Z23msrmnA5jdGQMik/SmeySwSr6Pd
NgQPPxkldMObze+QlPcxHB+vuxbcEnMH2N6lHkJuAWpZpc9TRsOxY/SQTCv19Ux0
4ykWu7s7PE0NicImakqNLOrEq7H/nomhQ5ZbEgPF6e4dIoQkDAzO/qQBn9YHkqVX
AYstaCgukpIO18d30kV9InDD4F5I4FEktBwhjC4pBSXpU8RRgUxPdah7lswL7qhj
BcttvcxWEhdRM94FYy0NaDV8STjsBH1fme1nTngUqVp9elCQB2CK8xZEhU9svy4O
JHQI6MKx1/DGU+1HdCJZvkfS0W2YkKlhnV//H0/n3cptW5/5vsQGD5nm4IYjUZqC
4u79jAqBQybi3JJOwylWPRJUq2IFbtTQGI7FEPWq/Esv3If/MIOuhar7sFVilTuB
p1H3fhVSaK1JG5vBPnCDGCGBLa7IdSnJiiO4ahj9aG+BZelZuXJekYudIOk7MGeG
tF/bLqu6hge2eHjjxvdjqDDUETIOZKZp3UdV27aVQqFwM6pKEgh91Akiq5PkStqo
NT+eg/2+yk4c79cfgyxzsr6oKGvKGHCOUCUvSR2zTOQg2oNh/Qm2PFKGtsRHMQgr
QL7ooAJhT5mTZoGc4wl9yp4hG8jY2Cb/nUn9ga9IXUxBWnHhEIAz2CBzkGastFO7
65TnfG9nkuJgM9hIgTac6Qfmmz+O/P8W2DAdNwXSz/8S6FKi6YVVbm5GaK807tqN
GpYkb2uFk9/5XjFgtAe7OMvIlWoC637KyhJwieNHJM5WJmI6ah3te+24JFszfmPs
50dP3QiogstK6yjJtyIypwZl6DJ9LOI4gJ+ZzUt5EXoQgEaCSy0skn5oePbgoKHB
CBCcbxyocPWZ7gJqiaLrNJVn/79ei1ET7fNEGuMxVTP6+Zgswxdu0ixVPuB8sMUg
YlGC9zffBNMxSnn8BRsauigtB2CEr2/w/FhQC45oK38iFqu2fsdxSwlUghPpXemY
g7hDxa+wet5tek1Qc7ZJT0wDwPArRM2GK7eyL5UC63njMg//TzmTRp3DyRTdcfoH
XhCoWpFiPTca74WDAzTrpo3QZpA2ABm17bAEQk6c+hPmdkWU1wcmpPiUpVTLTWBZ
bAMwqX+hyswd5sSa3hEg3qkwx7BleaT7A9aLeWhH8jFwjz42NrLgLXOwdcEa8NFK
fwJ6IuZ2NYLLi0TnwfjTRlctRYV/46XogW0pVcFg+aJk6kf10My0bVywNvJ7u54e
XXeTy50imH822PYrBKsHryFDlRYLbcXyvn+KsoQqrZOW+NsadQW31UMtPA+pyjkp
lh0umLmDQ/x9VqN3l0w5DMSBjw5oRbRSgNXYd4ZeVemT4H6rrSqttxqbGr77i6ns
zDwrU3atRNt1SOT2YkwvNw2t1DlYzzWB9itLrfnyYehpPSeZUQx71UaVzrYHnxLR
0lZSKfopxH8RBtZUm08WNwUHGpqonZ9GNNOMGpLL+qioVIo5SZiIoOrCaeWH3OKx
zKesG7zIN9hmQGHwNo91pvEmW+5kDrDRCw7PLWo6XW8PRNf8IdQKUWNLPODOG0PO
2Vh2qXsoohcdnS3MVnXaiZ7R9snfzwhSlK2WESCSMrfOndsjci577ZR77CsydCUz
JuSAJM+mbLYo8WNe07akBdmgrZ1AlcQxV4+ohtnrz0aTXBk/cNYJV9q/qmaW0Xks
mHOjMdaNdyq0g2ewo1qew1hL3ffR9NDJ6MuMUypCkECHs9zcuvDss1vueQdtA1jP
7Ez4rGWtSdoAv/cGJYUxvrVmSD9yB7e53HOsa13pt1wof3e1d72WMD92JLZq50z+
c4YCriu7qwSCNMC5Y+F0lwdUycVOEGkjROxlxrrC44Ay0eeMMlkSfFhfYgMoEhBU
9iO6vl0zlTC1H818lKnd5Izo2UP/hUS3C/lCpbcbFiZnHQp8l6MJGsC6wUMMj0Oq
2iqRXPKLjU5q9LoiN87i87ZQOT5nObsjRLCUXMR8ZAAss7UI4Q8wjm2c5AnznulC
mHSjFs4xRzNV0BDQJ2hrAQUL5hDP/qmNP2uSlTM39zxDNeGp6EUuzgyUuK7YDire
204EQDc8A4LPSS9Vty+A63jfuqrURPPcSK+zzzqBxdvhHX5tUHAF2c9+prLFrYHC
fsJcvX6o2iF6Be0rmIdLxA7k2GaAZWvE3tEpM2GXh3qFzY4qh0J/BbYRCHWOETfS
XgcLrP+J5k5Of/xXCLb+TA5YM7c4GZvwxSlGsm67q2eGd3OzpOgVtbkpAMRLhkM1
rGmzzvXOyzriC6mHJMJo32Lncd5UWv1sjwK7hHjzntTm/yKtC4WJl/7We4vxRHzD
v4hT+QOKqccS+GhWyJKa8rVUctaYE+7h6Q2AAxG70NvhIfuNCeQYW0rU1rVNL8Q7
6SKyy1SiF+zO1N2z43T9M9L3fqJQkUV5fTru2pNpY0aekfy7Ci/4pzHPw4DRk43l
jS7IInuBTzLQUFX0AYgnN/fxU9XfZYo5bjhEZDIE61dR+ka0AbuZ+xe0l9gOF0RM
DzSueAxaVZJL+p/MlKi4b47NabTfipDyNwwyYc4oQY1UX3ZFplaBVTsSZCfzfaz8
8cldw/q7WZfBJfDFrxsGaJpH9rIEt9mTqp8FCjRBjwc3n9afbu3PRFgaC88jW9s2
4jSGRyS47Gq1Cg/ChHwe62GQR2cB0Pupd8unCYm2HFzMmop9GnG0XjW7GiSPL0F8
wHl0+sF08mCMyxwGaCcc27YB19h4pR004+mxnOe6aKQur5yw14FvmPcxlqRn1Wqo
31CHXio2EW9sAqnumjaCX5v+5PglmJZJgRAS6H62L9GNOkeEVqa1LK/N42LT9Stq
qi/XnrInWMpBwk641CV1cCzTXHSDLTNVj0rdOroNHJmZE0d1/GeGg9APmA8j1jfo
epVJsseikh0L4g3qxDDGKQENZQIHmCoKG2QrvudL6ZJyjlVZTi3fTXmGHieSw2QI
nmsTcXAsHCUQizgQW7dSesohCjp0c5nkgE+e3Pdw/M/8KVbkBBjFj77qKiq5zum5
tmAQMNKMLaZqEATLx3tmv1Rx3a1OjPuehHkMXBAH3+hjz7tF9onr2VvrKHqj4pHm
zKTp5ISeh7cEn/TK+gZ5gcCAt0a0LgxusrgACvDhtpEsbzwW0h3tkLlM8+EOI28J
q2GfMml/f0cu8oQQMRa9IQloK2TIC8EGnaAxAp6kfCb9Oper4tOA5YmSP1yNOY8R
lTldYUzgQHjozukimhwtrYOJRx3lcE+UMkBYl3sfQiz35nPo2Cf1niFmepijHKAS
Z2y98PdvyI2w9iw9x9ySPBbHJipCsXpP+85mszfCDSJUBLb2PmzjEe6YRt3gt/da
7Q1tOYsqqOvisRDP/55bDICo3CCGCPGwiws5uT4y5/lANzpHsWZOMp3bHEMS8y1D
YLsCVUqPCe6ptPOdKAaidr3rarV4guzePoJIDy6LVupceb/4ZMb23uHWik+A3uWR
zAudGbx1Y7qn7hj+cLEFRy5EgYfon0fR95FaK84renkh2zvjPHeP17SyaVaDqv3n
TZbQeQ7YKWLzl0abApNJdFCzSfxbgEFtoAkQxZbN1JVO9M1oldn/zcXgHwzaIRMN
SSPct+O0OK3F4qkgo6t24rINEzcA0EJQydEoDrMmpo7WEkOmEFV8meyC1OCSUVe0
0PA86I2wmsGYSDMul1RhstFEUv2Bu6JVOvGu0S/oGVqGYXVOfQ6nHb7JMmktl+53
XFByVqFOURq+JYP2IyLzNcSD7jcRBklFV7GcYKnYsIYV1e9iJsmaHWtYA4Gfojt6
sgw1N9UGSP+8ybFIUsANcd42B6sdvJAXGA7sgYo4PPXHKRNTVfsfcIJwoh36XFFL
WvT+lf3lK8Vfy7k3nwfi9M2Z8JulmbB6bREMeeP1akwkOeyhgwBrQBP6ihoIpUYR
g11pQqw1QmydCDvZ5tcNrpV917YFx8c5hY4e5mxC55tlvz9ZQ2Upc37NY6bBAFzE
HDQUbcQdB60vaVS3BXR/MiJYf0+Si1e6iAiINdTyGho6dIgFb9gPckb5Nb4a7Cdc
YlPJUlkxivry4JbcwQXiDlWYwsoM/6rrRz2uywwQRsDDRwfWdXqIvbPbNvAY0f4I
gg7QoTuY81sQyo8drFwdY9scPjlYYaVfDD6AT6EhX/hzUibSBiV8HQ09pM4WV6YQ
Ctdby1wpIJLEbInrEZMVwKYvh2y/3UWVEYvn1vDDd8PNY/uinzrzDXU8SFalRTMs
klRnbPj6nc4N0MjG0rRJJ+UAfT0XMktutMYZYOlpxdLN2n6U8yH1emNg+8k8wH2O
M/dlu9m9GBmWOYn8/53uyPaqIcfqjhE3RegOqNnRb2PZq/As5sdBnjYRCxKWTz1v
JFH61eNpQodvE1zejGAYps81ixuejGU413/nqE8bK/4N4RTyxVhv5TAvKq3etkBs
AFzMZtNVbjEUuRu91h3Rp2tVCQLO8y2EfVuX4VLELTCulG6CpZpkxqMZ5zwBXvgd
Ea2fdIKUxtR+/QnQqPsnkEoD7jR5B8HC3UvASxNsrs6Mjknq+YaQ2vHx4ThcYTeJ
+1Vx/QEwr86AGG6NRpcvjXl0KN5ZmIGG+gWqwFigyV67UoU0EHGik2Tw7QA87/Qv
osf7yStogOvtiR9NUyTga+3DVqWXRWhyfR8joGsqsEuxTSCFomW9kEisW8zTF65Z
of9vmhiOgmLTfnTtAN3Hsa6wMlf+89SLantDOF5aoeyOsDdO8O3Qqm+at+DI0Mke
VzWHWJyezawuziYNHs4fpsGIkQwT+mgp8R4X3Pphcs6tSEOsuvC/2gNnMs5tDPpq
5y7/1XAeIn9fsDyJYZikM6DpvWmHUBd68T0uyme8pjapoBIueX0xLb5JpcjFbv6g
y1/Yl9cfErdQ/GvfW87EbUITsvK/s5IzD9pD0ML1/nvDghwjKFU8EEbjNDsAYdlM
ytQ+DJSP+t/B5lrYnMSIK76V9hRv5bL7RUeZkZFTqTJ/kwAfYyehXZhpanXErRFK
uCfYulBqXj5aFtPdOkI7RVNp8LcP857qfhwNJzwwzllrC+hVABJu+o8GSnEGw2q4
usbPbn0n88b1bvc1nQKsGJgkIcM2AdnCZsu5NhmliJpLbaChVIQ2xeozzdV12Ro/
sPMIn03EKmPDTi8Oub1zLv1rvrrJkxFay0jM25zEHDSBaXzaRTijwALh7SkKimRg
hrOP7LFUSRBvdf+LIQ2zQYaUG5HmHEwdhxBmfEa+KUMOrVdVEptRJJo+G5jVTNx+
3DWBgcsKbXT63wU7N0WZVbjJvUEva7AuXMRvT3yYUGJwh8AdjNRElS9EYfVfL1QB
nweJ4qy4FGoJQtUrPPFJoTt6BzvVf1JDsA/fXwnGHnJmlLEMrupa0CP/iFkdE/1C
kMfpHuFym6+VFT1mSaoAs9cQ7BNrujfdyPAP6jq9qmnA/DB2x7ZkTRXVqger/LLD
fKUqTr9fSAAU2erhqFCEqj2GE2twBI1tHoGbQAJ+AIuwNtE3jPguXgxet08jyuND
UZqB9WwIy8lL7rz7dCIlgPY/IKczUnpVupGvsJ65uxgdg2w6c2o5c5L7cWR9AtWB
sPXqH0booisP6qrcxhiWrqZlZ+fIIIK6G3Xfc+pHO+m77K3+gjPfnKHC/K02m0s6
PS5PhB5mCGm0FSjjhiqWEzcsFh6WeCymrOFR76XWsiWX4Jd8N++ofb0/V1hmU8Gd
odzsiNjgzck3HFu4t00JOlCTEbBMp2N1PjUvWCru20c0hODJ6Ym06Jsg+klLUJSW
NwZ/iY89YwGdKszs+ONsdOGsbDX4UNOmgaLIKZteo3WQCo6ajlrlsr2GnPzevOHA
Su/dnLYAlP8k1ptkiiChIZSfXqLT3XkOa07LAhmi4evlYXPjgeOkiGCiNJ8SblC6
4krdCGA8IB0LCu8yCJjGjPHsIAVEbiznibmLE3vqjyVfOYRnV78pnw900gPl+kWu
nm+pXx9vxybJyvj6DPp/7RgoefwEITfDkl6H0lcK2R4xlPtEA3rGJuxCfl5amhSV
UHeC+GiLxfSRkDHwD5ZKYilIDwZcAIxEwnajR2G++5J+CGZEQm89s57KWNbWiwPB
iWjtvzBlFKtwYGJgKxtNOPPcAh00A+d7/kx3j/955F1NL6PtDU2DD2OLkDzIrHX9
hnh6wwtA6eh1Y2MVAbzJ9u3lvQ6qFmpJno9dN0poMPHzIvqlPfjd5GD+lcbbZiaa
a5GWqw7w8aO0NcXKh/F+LCjmZ2J4OUTzGCLtnAK8G6XYoHuWXrEhR3GH1jp+ajn4
7blsJg7L+ic+H6FmmEH5zrZRIPqL7la8M0GFrbKpNLwehVh4/cJXkZsQWznjZ65Y
mqT8SFaPtzC+pM2niUFSLvgH+bLCj9pT9WfYknzOpj+Tmzq9aJpDlyzG6fw7eyw8
e7gjlN1zcMeaAOpcW1AO9DlKDJ1zLMJBNWmYeRYsUKJuOuvBwhi8jigHg+WB2rYu
1+kYUiyLLM9Z44l7u/1xV3QA9XCGNs/naLYL6nrF9pOrjgF+HpZtHFpLtzdiEZ/n
zuFvt/ADaGZ+4xqQQGVFK1IluuBCyXo8jKw6gOUbMHRW9cgZiM7JPdNCMRNjOL9u
i35IGSlXfKYBvEosIGM3AsOM1hZH5Ak+2wQBYB/UFRR6FyYJjAhV/nENXuF0BNnu
AdX3Y0TKkoou0iPYiYzJ0Eydo/dPqnbmavmLDPnTw3JkWmzvYIUAu0kcmz96GPf2
mBAsmlHJJBPWwUPIvoy6BMrBKZM3ke1vBCIZzmCR25ZvzPOrPv1j9Xr0RqheJ8GS
OtWkYbHOU7FIHdpKPYPMFGgxpSJ7+YEoypHAtBCxtisg0Juv+5P/wp4gLvVbl9aA
6ds9Ey4uoIuCJg725J569X4eMvCAkQo6NAp4CAQ/fgqF8L26OoKbzT+HvXz69kBw
1ezod9ypXKeHZHVSk2lBoLpZLwJSzw5dNfeDh1X2K65IUxHqEgwVhjDdDpRkYD8O
XoAWK/fWVh2TC6i4zyVYZjIChT5re8+EkJshOeva5BUsQruHWZQTgfrZ8QDnEYqx
f+cnss20YD8FsARzNgws7TfbCNVAZLObPv0KgYwE5waecHvNkOrvhng1bRqdRBmZ
KgsE3xkjrb1l+b0XO7fdlz6wYVPoN4rQcbcIwSMmz8omKJ9hhKuH01j8jOuWI2L6
zO8SpI6KN6Qr5bnTGS10zryVRM+5HUH0U6jvyjBCtOiO3EUceZ7RZFyUzEp/YXyp
6sfIzMDkcP45SHvyLJpz6XTtZMbCJWTmlQuG1aRA7u7nq16bJ0q67QM/KOgplQJ2
2J1QR9Q+zQkmRMPNNJzxfiJzBBgets0zm7XTOKYtKGOoSIXzCQYQL6iQVGFmHE9t
vYwmL9gRjEXGzmL309I6FrFG2xSAYPahJep7km4WQSH9BJocmuxHPNLei6Jt6OCg
9Rafks2jHOJifdeoRCF5FmFv5/79Xt9P9TgdvYwpTp9QJxZAYf8y4B2zJmMMgyeR
bKUaH5ZcXIQSyIcFrQAyFweIa5stbkXfUB6Mv40heowgUvMfK2Bs9+wY7zlyswYW
52Rj0lzYbLKl4T264KiNvscG/kRGjn3HiVeXGuTUJEM+4N7h+6iQW6W/d0Lue5pm
Oi0AbwOrG4UczLO+6v78/IcNvaRKF2lnf9CG8JZGTGnKVAEqYNO+3Rf4x3HUIJ6v
8Cw+/qd8hMxLn6nRrRmAxgBljPWprC1beZKdnpaXgNZhAkMkNQ3khpTxCikrsZD5
5edpxd6kqqX6pX1J/VOggFgvHCMMLgExP5DllM0ogh1U/c2PNBHETyXXIKwquc9H
lAMIgL6gBWIW1w2i/WeI/xUzbJNrQQTPnFLK1cUcLsh1iEbemZAFcbGh52CwasFL
Twd6tk5ryCDLxryPQEiECQzPXeJ94v13U6fSDPjaRHhee5kZvxUpW5iebUXykNl8
wyc/6erUYjv5Qr/o77k/o4MOhnBSxFWe8fxvIqyzQCn7a6xRQ1XYbUbQ8jTDLJYR
A/VNhYW7c5d+NoS90WBOUeX/MCFUgdNnUzbMn0oRmGdNU/K15KSykhzrLnJ7xB9S
0fb8HrD/N9Cq9Ri+N1Bo10uDO/yeCxQDGvM2lSJVRu6imE9O+j0eMJVI2roIdAd3
q1kxrWX8hBaSP4xTVGcOUuAkAbcf6pilgpZgxDYD9fLoFs3/Xdf/Kzvi9qbFZ9Nw
VvLHECn3G2gy52KXDj7vPVE3wB+Yyl6UWiiYDKgSN3fZgHGzKDtaLeDUDYeqTHVU
nAs3YJhGKvCC1jy9auerUAMKj6yh6j1ROGqWv3Zbbuwi7bhG0V9aCHrjykvE8hf/
3hG8cj9S611PEBAw8vgN2cFeCowrViH2XP6KHzaI5YfRgQOSkiOoZZTzGnQB9F8w
umhGiVUQLd5k3gArQNLyN8+LttA2BVUEsFq2pEl4CYrOQrrnXKMxaXm1bjS5HZlP
UexBoZ6zsf5zqP73Y+FRodajMXa2kGmQxFAf0Pa7AHa6sKIq+g4PG5OZcSita0nT
SEkl7FKF+X/PqKQ0tzBpqA/PNBdXWvV1M4hbXd0hrOCqqEwlOeR09KnivmuE//Jg
DtZhMm0gVTEaf4edEvJfeUgMW78vdDA2HxOIMHl35SaaEwXmK8tghBN8lfrWLGX3
BRVS+zGbWafxRDohLhF4nTAjcaWcAIe45VS9DTGNL/ziOlTKbSPGwh0iwsebPRkY
QqdYsvIn+rl1124D5LEScOy3lHfJnZ2mWsQIEbDXP8jLXFrGYXLFozPL8ZV7moNN
m6UuuTlHXOypBVpLGPGy34mCXxfwUn7oaMVfWw0DiUOXBPosxgEYDacstlY1FiPK
mo+1tdl5yMeGEgndXERWTfFj/6XDXAznIBEHF9+sEeSweJoGFhKBDZtEULjdmu5E
NCbvmsfYDMQqIy+/1CW9l2E42GvRgkSBR+X7soaIA0b9S3vEeyEdHNHprttDZyib
aK0QOx0CYT+DeamboKtTyKUWjGCuJoejuzFzsEp4/ESs4qhLxQ48YbFRTyu7x9Qd
TrL3HaCjePiOKSMD/svnmyGa7P/x/wjpHMfkBVMLEZFpsWVtWK+k9JN71kvuoHvf
Jl4ExXY3DL2eqmZb0KPwGLy5TCby8YV0o8/76LBFEPzNLMrrKS2MoTi6uHySFM7S
p1SzRq9+DovQjeTg0zzJL/0HaYC1MBjdEHZBGWyedr8L8ziRftTQCmXDjFBTZfNI
okZLaVNB1xpw0wvfwdmpag86XxPUaMoZ/qO53U/BaoKqCRKcAXuJ2H6+7hAnTRZ4
sM7XmOagvbGWVi2BvQivagQVIAZbZFks5H5I7SKCgakyO9rcNcuk66+Fcvl7G4dp
N6hsbRMR7+iQPVayMC1LnT4M5th8TN7EdXqLSpq1qSRmIKLN8VNmsllrw7tCF1ng
foKnJDCKBl37yQfltI8ZdIDS99EsIIljR9TuSSxD8+nATARIjeh3DWjqeGPgWnUh
ntcz5Xwf4e0Mwcjp2qrAk9zbS4Q9iO+cX3eKtx4caKCUBCeFyaJVSS5CaN2zXi1R
alnCtedDbawkDXUnMq9rtjP+jrLOizQYwkUUXxM2EnUMI6r2b4J0f3Qe4YbHX+r7
FHavzXpzf+17/yD/waD3dqqVLbL2ODqQ1lgvAAHB/sric1dTtGFYOhNcaSxybhHS
bL3h4sMQKwicESBHLCKatGo/J2yKm4h2jb8hkO7CGCcsFwxezexIuL4hv82EKzbG
o3/Tf4ucnI3DjaTKDPsYVK8VyTHcl4HpmbQl4NVmRmG6gVu5/fxZeZOD1bTa2w5t
+Q8N48Byg0VxxRZ7Pat0qze7FREo3zsqFvReOknZSe2llMwbD06Z/cFqPTIFacoO
WFbHebdkmZKk1+xLpaQXe6v/ptsGNXqyNZ8BoUpazGzkAPKe4ZYN/EX8daLj+cmY
+AdH9IbaoW3Vd9AeQD3T6QU/vRuNA5ohiy7FAg+G1/UXkryb4gHFrDgZ2vVRuxHg
j4aym2tKXKk3tQfSPt+YGpCQy2afxD1TBNYTvU2c1CIbNcHX3DMOzcMa34PDMEcr
LGj4S5io6EcptcknFd8girJNEzme95jaGkNMtzYF/Ut4Hmh+coX5wrsChzTJh6jn
/xfqfTn+FcUYxVd1BZavzsHewXhEQuSPp4VSOV/LSEN5Ddqo664PC+KouWw2TQgt
xCkb9Drk4Ab84JxK3F3OvD5GjgDvwpwe1mKjFjf41E6HtVO9ko2ZpaIiD89OmWFq
mgk1CiMt7dgmS7I5/GV+8XMNqczVHEEiWMxuHFabbBl78+5pDNacH0xIJwy6tk58
OvPiGVkFeGOWaY96Vj2FP1K1tUNcqkR57m08yT/1RHQ8s85sTbB+hXBGNdD0MnoM
a/FymYH4dkObM+lrrwl00h6dNaHZHEfVO0TCPStXG4DGmCw8DEbv4s1RvP0M8f/J
zwGm4W5OX/q4bijWlulfQ3nTnELlXbTHkdgveJB6LSGVl0XDbamLlZcmujh/En+D
O6hGm4l+GFzHpgUbqLLbANR0/3/U9gHRS5eNp8jvtt3/wjAJ0sC0uKLR1hoMG2N8
zfAu6EqhylgWsSJiMY/VGSsNE/2HMGML+stzbqBsz5BosaQ3MHFr/8m3pmAPk6LF
PJKVt4ktbJFRGDJnkOLrBbUOaENfUn6N3LAtRInT1kAoOn40CLo5OQ1aqYIzYXyB
ZJUxZ5qrodypKofsHtvDKKZ4U9fo64RWB9GvVjsmympLbxXewtpALwI8gvyldo8v
Uph2EPTqltTyS6RTXSJeyWuo6VfoBaGcPqygUh307pUJzZ4DmMusVxHTWnNyG9nc
Xy2LYWv8mtKIGWdyRJZEG4Gn9UAweV6UGIFL9UYZmkkzujBt4JRHIgTNZ8OeXKHA
gFnomn5QWK4KUoGfsI+9wf3sSxRzpCH0Sbefbg3uyQyO0T97liFtlsvyURWxmgbo
jbVq+Rd1AmzW1MfpcQzju9xv6U0mDF2Sbw0l9UyPs29uvJHJ5KM4sfvv1h6BVylI
cjiyF3mVQNUGS9jDcbP+htOfwjZVfW9rcusu+MKRs7qtI+AJWiM7PI30KgMUhLl4
iuQFp+vhT0ML/xdC9OwPJsnEPXBMfNPa7y4lRDInoPOA4DY96/xfDibzI0L7iITO
+G9mebhGt/20GxbyXKr2/MSWwB6iZZxT0B46LbC6wFF3/Wt/lHrPvrWRPspkTB9H
0eBc4utDHxY4wXlGIAQ/3/3it4nD/5WWRglYVO6VKEl8AhBRwF1d+kBdwSl6imK8
CORzlQGqrV+3LjtzIqsZUmkw8dEEpyaUwjqjT4zIX/e2rACk9SmqwN+5dIB+3703
MMhbilahlZYiW45UXXYLo0/9z+/ww/CxWfGxVq9PM633dCJU3cSma3Jve/dm+XiB
orbiUsHff7gIekcsep3af4RfW+rfyqCwVH4kkrbd/ApsH5ecPOw8DfhazaumlEXt
ms/3lp3ul4Z3h2bR/dcQBOZLXXJS3wBgJNIA9GZ3+r4YtM773K6VNRcrxlrBvMSi
dQaYI6B6Xgo0JrCAnuIZLBUP3NiuJho2H6SfySFFK0b4HNSJW1wEb3CPEJC2+gi3
ha3YmgC0MvJ0X5Wq9HCmbQ0q+LiR19TJG2C6hGgRTVvlBRBJ1g/1ioaR/fjebqaV
r+6707F/2et+z2HVt9IbAii7KqMc3zRyKh08OQggrU8RXfd0JPqH87Ym43jTzb71
7uQu56kUPfmn1J2ymQJgtJaFACMMFd5Uh/VQA+9uLtzT4zKpw8tXkTaXNpr5mYCJ
N5/dFR5DgfCnT7tAMvjFHr6kxM3Idmwcdzo05Fr3Wa6Hn6rSt3bgQmx/zbvRk5ML
zXngVe0EO5Znzi+PSGOXDEelEMOZ3PiyDI7lTdajmIlwuu4NX6R4Y6/2iPugiJlI
r+hdmQkFK39nyQCpUBP+qhpey//W+lYRtCh+bjiBY3zjUMqnxmUvHJcCJ1oN2rgS
LZHTmQhQageQ2+yIrFZtOwaDYUKZmz/eHKts6z+Akps2E/3GwN0EKSu0FiJS/Z9g
7VVoUjdfWgs9samQa3VF8xr1IGf3GHuxqNpODa0uocMI+WVY24BS/+NQlf/TeuMu
a7rwTNDFnyn9Y2UTkCkB1E6FjgRYV+lquwRXFVwI7TgMBqsXmhDcRZq0uIitcmJ0
w95Wfh+tDmGzB5AZo3OvGQK0i/wP/YZmGJypXMUMA8NxyNrqa9xeDNeWcV01x6Qk
ZfjZUWXJj2u+R81kOjGMV9tf5MAmKi9dqa2EbGzArALcGexmysVhF/Di6CeiIJJ5
/kcYRd4eB8Ui4pvpKwsA/AtuzqO+bJxAyb75M+b8b9UFb8kvOWHcUV7IW9ycZw1D
ECpeXztBuBOdGIt5H4Qx+anneN2WsfJbGJmecxxP5NCsbXwWsPLDeO8TCfpf4KOz
31X0siTuBKnCi3RPDW8SmAOwllD4hsc3aoizYtLwH+o8PG6ThJ1atFprW7lnl4ba
VE7EGrqQJkkznPys8K9WvAQ2pQYcWj69FzZsI8wZv8dwf0H7a8KnYk+KhUPRFZyz
9XZDpi3gus2EtOCojJNtTJ87GQC/ikmJlF26M2fmrmCKk+L4+xn664sg/R++6p93
L2SbFZtYCvKb7WMBvP9+iEDJHTcDjpldzXf7v96/NY09QSF6Fp+eETh7CM8/qv1K
73guQYVNHsh+go2eYs+d5U8odXaBnMVJIXdIWkJWkK0SHsqpX7H6cscznKjqPEIQ
lxnP70tHPUMnJa+KEpsXdQuDpUR/mF5AJfH03uj3V4zk6a5fGBs+TjymLuMlgBLd
0Ojr0k730ZIq8MIjqnZCpjDJM9wMH7FPKWn9rOdH3TMlBUzol7oOPrkwi5goxon7
FBq5w9cfCOl1fKSKmDQm4hCss+yF7ohJj0LYd2fabl3ZUEuM/tJ+Yqin1MShYmQM
lru2n+DAJZDrrmtp7MriPkz8vyzgBNJ9qZfRYGsB0FAgPMcq1G2rTLK3bR5sCAzv
iT1Tc/WS8QNddsATFQ9F5Jcg0tehr1y1VB9RELx4TtiPmKaM40zhqYoohHG+LwDc
miHRuf+jLjI7wwsCiqatvO7egNVLJl4di4jfmaTagOJVKhbbUdyuHNUgA6wFIGH0
2mdyxHxJczM15HckmfiAx6s3DUUTiza81oGMzFhfKJHyh4n7MFTY26zXIv7p3CnZ
VqA4/ClceCFz2Dsh1GTCcIyKDTVGwN/kKu3I4RolciOZRAIIivblFCRzIP/IShwL
A++dLmJx8vygdUpQUDNU4WGH13MPg0gl6IdAqL+dthjQAyS3Z+lV0S4+0yxrvXKZ
znHekOh5ST1hPHTmPtulSs1872QeeqSZhb2FaIvVq7KmQqqSTHVM41xKVhgaeMGu
kkp2Yq5fILaqfcia71G6y1hcrIBh4OE0kY1VsvMyzAlnlqMxc76EuLLyQUxZ9DAh
la712ozHfbAg6ePtHLD73oPFXVK6D7HGxbRP4CxgqLS6QwJ0mHRm73WSfuVTWbXZ
6+kfWyz0OXO0ur9nRERaAOYu86mE78hZl54fmbVsXO9kkFZ9RWtWKJen4l5l8xF6
YNqvxrjwIFVavWVBXTq0CU3aEoG2jLNLayCtdHL3cwR2DO6a0gdAspUQn+6Ce7fB
pDJRqPh2OlZky3iTipS9/HkTSvQuPX+eJsfNzB4YUxQ8wdpTG5nSOb2Yb5i8fMOK
EehK7hQrZojT4t4EftNoIVns4Fw0BrbSl/cNUGBJBoITLPyuuKH/N86dnKb5+tTW
cCpb/IFnF+9qC+cRgxIACVjzulNh6P346TJ8QJur0mfF1jNaCHx+ACNDXOt3OO+E
Eab1XH7ud5Jkc2raP+7udobc12ptOw8/StFfZheJ5YavCzlfi/3TnbAaz06ik9TD
Eme/LxKLM19mTW3XA3SSqoXY8M4oni9RC5urg/ymh/0E+nasCu1Eb5QwxTRs+znl
M5nYFpWHMKf/w+CfFvhlwYOE8sS4wRDXPKDII84+Ivywwp/0q25SB24E77EKJ1vT
O1I2pWiHSKhJAaf2b1PFEzPj/0c5QX+XWjBXqx0OMGubHMquRCBayikpw2dOlqeh
nd+vNIVkDxHrCs2NerW4TyCK+y3Flvg1LelnRJTwo5lCTv2uDXi0c8P01RB+LHFR
qU04+DBAi7as88ftPWDekrZZiNhlKR/ie/CGjcVzmzYThqjDLvT4ICwp8chdnUdr
r3WpW6lt8kkQWBQpxX1Ohqns7NxDhqUqtR229p1r1YcmImzzE3DBLMIYFgGzX3mw
9kZdqCxLqcB+bdyawPVOT7k90V22NanM9X1tJ56l5aVjrCwQTTLfwV5cvC4erIom
/cgIS6hGtkAv9nhTSo3F+mJ3F5AzCHK6DWyrvkTm1UbzeKvALSP+QlH513w7YCZR
MguyURmtWkGocP42mMtr5Ii+P2TwFgVMpvJp7WQ3UYR+5uX41PZlDukAIcaONpCx
7qSIX/sT1ff2U+Pu1qCxU5ffpRIovKNfWH2I7HftVdfuxeK3ffgae8tPntl0VIH0
Q00XV1MNeaKnPzQmjssYM6WLOqNZQ9JRiNHm5eXctgDm1oL7UgEKqUMAXv0VmGcZ
mFx8NnxMJ1V397P8VISnGJeTJg3ScmhzarO/N1zt8BzTfmls46WQfJV51q4Jc19I
6bG6GsWVEdMBGxz9mMhQbnsF4SMX7DVJZPLrmaGTlBq0scWrBB8kVjrz3gbGaWPQ
tA40ylEGqU+M81nBAMWOuogSswfu8ji15kFPUoT/HcteNq/ggOwx+U2OCtVEnNM/
3kFx7wLJsfJ1567kRaCC1AEaTizoBRR3UMBKDVyWBVuGEhex9CP7wHDjV3sxa27Y
XJ5yiQnu5BBEYtWHFQLmSAwb8u4f52gzIO6bEICoUVlYwJfxqu4BBytnbIDDNuVp
FzKJjFvplUIlIwVC9VJx1MTx4Flztq38xetSEMYXSPZI6i3QggibKnSkomARiumM
AhNXcFkAuv90FUXb/F64Xy+P47sQbreA/s+HiiaP5A85YLkTI9wBIdk7uJ5i8Ma3
0mgwtgIo/GnQySF0xh8opNZbQ3BGrxhXK75R8kvRNzdHTh80xp6ujKUCqZVMFwx4
IZx0WFUaBC+3BBmJqQ+eXKWAtM6nPrTfGtbAm/PfoUqg5qOFawa37ahIA1IxgQTX
Bw9dHAbyjjBINsQcGtCSqtRxq6XtLCMq1iEr4FbMw2zKbZZPFNXDffANJZ7eevsA
qsDZLr4CumZMfy1UJiSyBrvh8IIGZAiJrP9dseyMVtH30pEDur6jmSXrUYXbQ5H5
AIfM/o9f2MlNxoc3AEi+QWPFdUqqxKOi4M3HF+jD6CKWJMYME1f/2zkjjKo9hcGb
sizgaE6zLVam+0IybQkk6EBcYhIOcxufgr98bER7yWEvwtQY4aS670YDhBrw3ysn
Go+cMc/PnVln0lw4IdwChFlukNV4o4u4r7OGnYELVBV3EhdHD2vaZlcEuGGAg05M
VBC8nAhdL1aY3vBa4Yy9zLUV9H2zXP2pxDfZ/+7UZb3d86D/QFY53JxTiZJOZQaJ
is1fOFGKmwxClcIIuDFNnW1Aksb8RTFzlefIDAJxb1x9+kPi3q8nglbCpT7bh+xj
ELihljlG8aID4xOqnArbK2V/X0eFvMzAbV9MIvauIgvQLGvFToSkG1d3K5JeNRqR
Z1w1XfpzLDToyKO0Tw4/jVwvYG5Wf0/NJbl986yQSrJYX1kDZhzzUdUBN1C70u0U
2Gtz1yVhCYYAeF7gwhsqBMK6+WTQFRyLfAq/FS7lWRdSIAsTG//+bmZ4HpkTlzvw
4AlMlNkjuwQrxxTxf7G/NKrOfP8kXNaDMLXxotDpeLL6m7tQW8qXNsgHVZaJPPL6
jJuUZFWPkLqWlUXK7mH6MMj0QyU76Z0zJ71rJStPoRLEr6C08Yr3ICOZ2n2o0x7d
TYL+O14XmVnSG3LmEqBqwGWC74Ur303zE46q/EhaF7/bwolmXhAxbcMgi3RHFAYl
j7cmjS6VAdRnize05SY9oGML2sF7rMxntiAftCiK0Ipz60cL32zzUmgZ7aHrfqKf
0KSUfjSKQ+PL4sQpLT7dexpzzFAHflrLWRRTGitmJbpPz1W61ZGlB1qVgwh/uTfY
dEQi7QeNjM549ABEIeFZPsVu7VUTJI0PsYI+freEQ+Y2x+pcGeUdeGchdnfD0nH2
e7lStJrDmPk5qTTIQv97Ml/2fI517jC2mfU3ffGKzyEKmzzTX1k3m0KIzDDKKruZ
3rVJ4I0uN8NVB1jcY0dTgL6wAy2bOS2q7+/52oyBMpHwOCaIwL9oHCAnvr4WO0hH
utF6GmdgPhqbLrAJn7nXf2gKWOClQtSYM5bYCyJdV1T7lLGuyksIm+Q66wuW2wUY
lE1DAynLNtwPNMwzCHMezlvDICLLqNQzYQskbuOYlxHib6kF6hLgORxk7f4GUAXs
AHOby3WpDSirXn913SRKyoWc4PMFnxAkNbBgd9+SNOI1tNk++dc3j4HMC7KNWzos
TxjB/+C0sM9ak8VNPN5pFiPr9VEWhkJCBv7zi7KLlSfi8MkQGFZSrCGfN4/7yHHI
SV7cle8brBTLa9Y07q8ALWSUeL3FSe7E5F+p9Xl4/4vlRIJ2NkP8DWgI10X0zQIA
Hl5mKeZPmxVjuZ3zf3qVyFd/EAof5zmdvgzp43u/i7cCs3FUPtb69bodakNndSf9
lTFY1jLO+O13b4cMjeVBE2qS2gvRbuMtZkSLFrkg7a4nJHPPDRZxIPvvst5cCCPA
QOc+slo1ykChMTdEXs5iwIT2KDbeRm+56HEeeYsimMtGD1Q1zfevBf+IA1ZopCvP
iezEUmV49odtN5uO/Nsfg4r1hZHYn7wyv+qxuK13FuEmNxGlRx01mlEffHjEDVZj
PJDkTzyLr7FkZ+j9x/t2ua/vay2+gSN3myOUpdkoy6kmB2ubMXqTvIrVVLvgCZ8x
Muwpk+fm7/8ffVCzoBwm40jHTLsRr7tgAGZ9xv1a9e3sXqg1PGd6uYXYYv1ChSnV
graN0tYNkP48V+FRQnyrwvkXi9efmg6ppmDm1gVxytMNO8WHeGOfH+aUvhmSB69M
vHrJzX4jXnX3I7mdBVgkQW0zoYQ4RQdNGK1AotlB1PzJaqdefqpJPuCVvUUQZimG
OtVlGGtKgUqGKNkj3Zw/rDMOjWZdmOMS0Fh5O0KVbflPAc6MaopfXj7dP9/vIoET
XcXGHTqDeAxS7TeVj9F+9DnrKbpJYlEWsXfxpmdUeYCar4tJiNjSqCZKnk7ALmUD
ETBWbtbYCT9BokeHL/dT3P4fWhgMYpubCMZl3d/zfukMJGt/6cyONUo1/FN93Pjh
JyftZu9ezX+yEzXceTKHP/Wdxp2u7ke7tMLTMrxKQn3/VcJvYZtis/REgGAn9+Pu
rI5bKnNFI1JuTuFmcX70gx98RZSnR7vaWBJoBWoi2FzBIbcJAhFmXLv+sgOqpSeH
pqIUItIG0yUTkLcUHEm5/+wvfSIG6/sYpeyysHMlmgZzzz+3OGcfIvOws8pRQrU5
w9GpuVQUxnP/wRDcCVpBCYecx0lFdop5Z+HgGb23aZMIktArtfx8nFUrOq2ZLPJ1
QuP5cggxjFx7E+D9GRMMs4nktFvFHVeflIeQDcmiVrLlJIGFIIB4HtN+W/C0DIs8
k3Tw21CX70j5ub1LHiTAi/AdNhuabd2EoAju8kx8AWlYTf3fA0PMnxh5mfgcC+IH
eji1w2P/5y9SGTnXR2ZAKhdOPH52KxxOQ2+v7B5TCjSlAgJofVhS6ZJtfpojp18X
GCbbEs7sgTy2VDxxAmTeLr/JKXnd6k6pUyeZdibAd9eWKnDYjYQjY6iM5rIm32jw
JVrt8IbCUQDlGEZOxAw/0mvLpS+jLF4Ge3n6NF7SCCrA69Hc7ccTmq3V5oPdmZZR
2KR6LXeWFp7ElDBCunez86KKEWZTjSW4RFFg/C1GPPobrOyfrpD+YPoM1mt/D1Br
2xFIreYo3PmSaU2EM0T275B2+kE0sjXnQsF5+tY6FbrdK0Ul1Gc/Hq++0rSYHmit
dkuGGOfDtw7kK8HTUccmVWhI4iRUYvgpax4V59V16YGq8Z18u/LCSkx+Azo466OR
6sJn2pWMz/gH7ShAeeylB0duXst8BKmIAPLaR/jxu9xt89KCJWIopx1zt86J3uPP
1y98tv2Nu5MwovIF9jhKB2NOOVbgB+TCncat+Z83YBgy6oEHv5ftjRvOISpYqoaZ
3R2wdBAVTivWHLutLFgE32T6xK9HuheI1inr6J755n4i1it7ossE6C+/3t6obQ6L
bs7MuaxGkA93sCPc1u3mOv0OZKcxxZUw2/alRzwcD3mUTNhTgACvRjQsLt5XcRta
87WhzmNW2PiwTpQ5/AkxIdMh2rLhEUWan1Aj/Fiy36+6kX1XLW96bClr47VKYt7K
JxRlnfSVbCcXSXvmkvzQXVNKlRCI/Wu92WqLR3XkTMMDKKElB9yp3TppoTLWbsIG
+S08+TGodXM0mrWbcQtZTV3L80IVl8rFPoXtDH38mN9Fto6VEqD+ejjoVI7U2ush
nIVri9xJ7p/ZK+7oHmPdRUmf2Ev3U7DsSPmFDyG3SwCBpqj8/2LJ5dK4GQeeDqcp
6RYKB9nhvod3donnM3j7ntQbFwf/7i1E9V1gxukuXGCaQ/7rb88ovBOz+b6Hsudx
xkc5Gga4OMi0THe7b6EHq2xbA79cgxO5jRBeG1/+2ihCaOoDEc2tyuckqUZEg80U
knVmZvRFR0gRXzEKH1/S7fbzZk6dY5GTI3f+DlSOtUrVNbvEvDb4v7aK2oK9VBaK
LEmUyIibKDXpCZGSDYIWVTI9vBg7wfeFIYAL9kCluOpyJFX1WXa68WL9JBrWOf07
eG9CXW7BVskfFvGQu7NxWZgRc4PvJWlm+Gu8eNVw27ttp9FGzK1Xa1GZ/0hzJUrV
rN1d1CssdzAh/VTQd53YqpGTRBzdsgXZhQR9vvrXWCocCA8OB77M3XWPZfoZfNtv
G2xJAVvmM+vMOz1diZuvqG5g7MZnpb90WwGU0AwXwt6cuuMRRNEM/A1GpWoZHmWN
WcsgKKQlWrx5vZfVAFbO28Qhgap1YNmUAtk82pzpA9CWKdVznCpL8FJFpEhUhT7w
MYqLMNE8jleWjQ90+I6TUoDchSbBSv0SZyUqDlzmY3823yftbD7RydSViHODxdE+
jvz2tfJ4p1iOL1GYKrz+XUcjQtUP8Wbp0rj47UcJHT/xD3ycRTd/u4T2C4C5I6++
+9FX2u/Jsfp2pYwrERXgGFbXSh32LbKqvFJgjTVxYQqFvyxzxzLkRHb3Lmc+n1W3
eIB5gXc9o2V7aMN8UjHC0bDYh/mIv9a3v/ByaWbXkdy9u2s7mIR/YXw1lwx+DBa0
NDvZQ/qc2ZoEjhhQILycMMYrrzEMZZ1Pgxn2Ihr4vhe1Z0nJoBbAn+lwbR95cGt8
hSY5s8sSjqni/6h6ONnQ4ZGcethSpZ9HM6g1JMMDzZPT51fe90z02DRfmi4gQt94
VMNCaIlIK8ABiV/h7hDzgUcdh2zrg6vPq/GhcTiddy7Bg+ZuYnWNCTj0cy6Ab0yx
GZhyvnb6n5g0TC62dEEG2jTGH667AGZRp3j3j27jRGV3O0ZRkaV4Zsv2WVnb9kkc
hbUAGZCOw4i12kMYa+Ryup3/+7NRyIL0pVvzimKfLKcI9TfKmdha/eMCJAVh+/VZ
tgrful8O6RITqNyI8wxe3fpvoKaTmToO/gRgFGM0PKNDVMfnciPAYIpLwbsV0VJi
J9sxwhR9Iy4JJRTCPGiywcpvjs7rLSzTaNHBr3RqCO/h6JNVgkFy6atSohMXLLC2
1Z/JtIGALOqgp7azS+AyYTGoerCv0ClrVOhqLPch4mzCJuJEUyVJtBow/YKe3Lc5
w0fPCUfz0n+1xvKJaDXFLFI9WZ/VjTwY4TS/3X+y9YplMgtYamFNU8TV9rMQU/IL
9DPIpD5x4ZWvFGVz5eNF8I1EmN9W/u3Dv9jHFP+RuAmT8DltqiNJsskg0z6kccpz
Cgd8TiK4rSx++yMrKdOzUAtcTetPfgNovfmskZj0XA5mgCA6LWHrvLTw3ZbkjgAJ
/qXfK3I8zHUAhSwtgYGGnIu33o9hDqcj0YkjzeFxoaQLmW9Oo7dQwK3rPRUyV+bc
87dDAHRD17f7vVHISxEDRI62j1snZrA7sSuQVE2fuaX0knv7AYx6qFDeUQBasYY5
VZNRiElGaKoOCeNPrFp8AFRZ+psi1h3wJGeV50InK6rTqcB6C4u2XF/GV3J15oqe
RKH+czRvK2e4nSuZosJNT01cxV0WWsDel0tufmHO5VgUi5B8WNAykqWmT6zG3Tsu
r/I3kU6BCqZUXd0e8DvKtJGKqC9dkTE0A07WIoCNHtOGSZTF+KV/c+Qnz8D1d+GG
IifgWimCdJe+cDVoPl7kaQdU973QLt8za7iDkctCd9+Xif5vmGguACy0xsYFlFfL
GZx8gqMOwKpQFkAQRWPd44e6aRYZERJb9z5imP/Ae9elYfeb/2576WgtbJ7MVoVu
TXj3KL0pECIeTPGTbJOgNkJd49sGPlYDLhCFstQRCAe0V9PhV1stqbJ0LP9DCr4U
H2kzXemgIM+kKUjwYQpaNKvKx6frI1tftOB3io85wTnsJxW3c/3EO+7vdlbaWg9s
NE+fCmMZIIe2tT0Kp/uYgtdjPxeDK6Bnmpj1uJCxxQAceZh29LlVDFBKSjnL54Vs
p+I2FDnPXovEcXYXPJFatL2hrRg8yVWeLmcieun3bWqpImXs/PTdCYuSFFA8FJT6
gpi3DPuADCh6aCL3Taj3EPdLmpzVwTvB7CG3WZU8x9eBWgsHOJ8LmVKftkuoUahQ
clVmhWDCjCsgGWZMkKwfNVwc55pGOmCH5YTK/qwdHmPQ82MuED9myI9SywyB5++/
SbgvxYQ6bJ8DhTBmplZxHSl4h5Qk5SHH17jNoXsD7JTWHnI3e1Pb6uyN9E4ht8UK
TgU/xzK0lYT5Njg/nd+IsBpBw+MM8beMd0rSNTVGHwGk8X6pHeDnKu6WZvA6DMP5
D1H1Iu32oge2HrjL1RH39HS5CDS0VH3G71R98a2PVk/ANMhR+t9DJSzkHCL+IMVP
QHgv+bMScX4V55KhH5I8BI1vF8MvT9yCOwywc/xAomI8YpcaKQBCX0H2UjgDmUMA
81iwAf0MiWFQEg0IkYVYTUJMznNtPCWLbPQ1gTw7NPBJe4ceXiUlr/DAYvifN5y0
1Jnd+3KSXSVGJKuW6JUY3e12REObFvIWFwjmvGM1CgO8UuguLHUPmP0zR2NyCkR1
kg29DLPIeIQ5ktDNv3zraR+wfou4ni7PFWz+nocus6syndqwzi/UGU/2npe5BtTi
wX2G6O8nNwO3gpWcz78HRvDp5dOXEoE5fTZPehHl0kkH+sS79kByz9tRD8IhltsR
HivgrBXO3stXVl/uGiuFGQ3+LlaXRGhB+//G3+ktbnsV2Zn9OiBq6O+fzqZV1iQy
NvKPRKBl3IeR/N0UknDsj8AzWZwef7UBsXUq3KZxb2lwFrTKe5Y7jmc640yHi3du
PlAsXJAKd9F9MR5H5tEijqJfztQd52qfyItODV/yjI3rp6zZ11GXdjBb8TLcVUzQ
J9fzgCxgju5z38Z81a2WzmV4wt7IFHDYrGg5dc1icQ7LPCdm8c6EVgjkZhLYsmYw
x2zX3m8KiSElTthqLvdkrmXVxLpFoOimgIKZqkIxEeRdZl/HEFSxZMTJPVvbOJ16
SGP9qcrOEgY89zxfO1FbSdZnMBm1psL6IcqowY0TLKAhcxOF1HbF2wDbwSQt9yzs
XFnty34n8rrwPPTFHmAcE4MhKDlfbABLg2cs/vFzVp96zKxsKYKalxcz8uX9wwoC
H8gPaW3Sldv59Te5iCpsRfUd26bdQfDtg3KCx3DgkDMsQwrNYoF/ENHBmAepJwUH
xrZj9GmkvTQQVb7a4sRPnsz6IHv46EufSVw7yx3Dkyu+j1P2WC0J8crK6ZfKp8dt
8TDahYSpB2V3YaTLG+Ze1TBN/G+sfy1E7xNcH1l063s/R6lD7fcVgrDGbobTCxw0
XPp+8kCAEPTwp0cgOCZnyt91Qk5unolaj4MPnDNgvNmWqwcv1/SVqoz3VszfPnBN
9AeWOamU010fowcHo5EBjo/Q469l2OxeSeUKl0dtBaaPSHbmFuiVhRJm72HO5pm5
PMqgcZP2ik27jMOwEzOFus1FD+ES/z77ZB9hs1CbU/HUmjfKxEuQ6VJTb7gjQ4GP
dEYWQ1fJN2o1a5Ti9K+fU7f+A1eRfXyMipTXpGQT03toWLjtQzYEgd+dHC0oYBn+
kY8aTY7UfN5gjN24mwB2J8sOtBUG4WIMMPhkdL0sJI4su0VSrswFHM94/8piY0aT
LJHTuvizBD5vR5+sACG7FAWtQpSPZwX2ntGmm9x9eeFaNdkgFF+Ns+gHgR/ouHCv
i4oebhC5rwCBtBrjpALq7rCwFexzIwDYiiPxYFYuMRl47YN2ofqUgFfIy3dT/opp
ziK7HhF5FS/ATl6MctFiddrGSiVD5YU1ohm98KVjIYHfPzNgCH0lIrURFATpUUTg
ZkTexK0v0pAn2Zd/43q5PmGv+eRG17DPrb1eIWGalbP5yw069VpDfJHvEfoLnqq7
hTmjpIthTzXh67RfSHy0Ts8U8y/46p/L/LDJ9Y1qPC1UUwrQB/g8NKa8ni9yXJwA
tbNSfrA2aZLsT1oIwPjQi4Kj2m4MochunxCfDkhoAZVo4SNNRKXlH9bxTFCydToe
XzXkSSjJ01sEM/aD3orWMwRrN+rX4h1JUtZPiU9RmwC6NdW2UrOg0i19ZNOo4YAZ
Y0UwPA1cEaM0mKr8TQrxqFqs2/skl9GXtcl89J59xTyFLKHZ72QJBwVfFCr8S4iy
YhUU9vK2AWxgd0mFQp6R+dk1KRxXhvwhXLdG2SsQvNxaNh+apRl1zBvXODshYXRx
PdmOrcFxEcN5mMySX370WyFNuYpVt61septCJlWVEm3/SmUp23MkIImKDE7juB4W
x2uclVtrZ6zNhEeCqQTBC9MA2J3YZqUhL2OkOzP2uW1hoKDPsfE5NDCkyg6AA445
iNWMVZYORc41JOI/3SbEU7ytG3DnQdwniKKF4EF4gnDV+dhmpboaYgW5Rdnqi0eV
m549y7Jb9pfBQIa2lBwVn0N/QQJjlCblckKS7P0v6kW93/yP1qfJPw79IayfeocV
sHCe5PACdcZQJMVpMMehc6UUFqpJXqi9MUFdt2kEvOPYbuxT6Z2EwIsBLGNHGqCc
M4DtLd+EGd1pfMBTUZxOnvMEM+OjX1Tt6FA2hHT1kf0yD55tJoRDhFXJkMEtYGvh
stfMlDaOGc43C4d4ParjghQ2x8dBAPZYBFT5y+xTdJlsc6/8S21i3mor0X0bA+TS
94dsFXTDEeihC2kn1PVBK9rXOZzIyAD4FIAy1ZuSWNg9D8nOLMszhHgZZ62Zpy6K
OScozgUKmdvkZIidYnzYFb8pmmDfSmU+JmsVnI6kZHBN4w2ZX7DXRKBqzLbhzwzB
vwrYqm/W4lgkSOW0Sq1HZeOkR55U6iM0GOJAeR8vVCTpRHl8+r/ES/D0dt3IeF7C
2sqemqBrZjCRuCVD3X12VkKRaGTql5jUYmVIrD6ZRm8N/UYBvCNuXW4/J0uSHrMS
ew+LsHqdevW+Xx0TwFdYIaeHupo/aP78715zbupK+EBwV+mT4oWAb3fUfxFMlR5v
PNXPNItp8yeoPF2gdsjCMr9FerNdw1yHQkQ8wYMo7zj7EhwicV4fX19ozAemMvnT
Swr2GWaNd+S8PF50TSao4FnDMvmXQ5Dy2Db+ZvwXHGJ54dQFH6VYUPi+04PfAGAy
OsWsWT7MOIuzSMwOwcqb4/+gdW5WC5EomqZZ1tvp4cO+rp+SMEYrFUYgyjkBsmke
mYBsJYwaP9ctf05LRodtNGc+A2ypsLJAblpMTovp5mpGNAgkB8esZJe+iAy2CKUd
crGdCq9B2AWwDCF22vGeaWz8yd42AKMveCvju3PVyaAgMl4FVkaNWQWqhgfozQxQ
Zrwa7xaxvJ66WJECCjpcVtbwUkV7W2NwLCiR0GFTZ3mzlAU5Ink4Tk9OSSpsbTK7
1hwaWGQ5bPF5IIKbgKde8GCPpqEaBOrj7KZ6NP055rYFQVhcWSGYtttczxbeGCxV
0+tzRjPE4Rv23z8sgfoBDl46OsS7bVX6eRIlLiUBs57VCaStT6bdfwKQFAA+dwaq
be8I0OZyPAVSRo6lVV9sXTMd9U3SdV3hazhrWAk4twqj5EXHFvOg+DCw9S7xm7YH
LZwoeLMOo131NVBJKmGfB0lO8XXj45xgjqcFwg4Umb+UJ/3fBUJXE6hpiNXIR40w
JyOqsaeZ1llHlJXOVLTdfhEaox841SGMICtMRsxBn/gxK4/PiwV9kVJ+OgnfG8D3
aiJQQxmuNM2On1wtx8ryS6tF+fUvaU+vk/Tf9DIAiEiA1tikuHPDCP1shSlcD6FI
hbinh/wf2KF/OBu8T9N4fKfDy+R+tTaNpVgZ2w7q14W4QErlo69+OM7z7eSbxPNJ
UwX8ydLGdBeDR4KDBdf1/HRKYZvXkoR71pwSdM/RUFTIBWfSNaxVv+g8wimE6ZZ4
dgnxtgrOQuJ0mZLKUXrvo+owKZGV30yV8XR+7bEPscJ8n+NsKIgCFEwyOKot0+Hh
PjBa/jrOpJt8sezRZEkMUadhg2jCCHWcO0xbtB05QwSuxyN0Rq1YueTXQi0Z7pVe
qO4d5ZuhQLmcULp45eGwy9XraX0inoAYlyL+BLAXGq/bb5pJ9mHRFXlzgjM7kBah
UG6iluAiEST2IQsQEEY1dRsqad/G/PjXHb774pB1BfBJsY9jrmxEqAd9zP2vRHz9
mbJQiuc623yeU2PdmTYDDPbucL2ziluuxreDlR2REe/CFZ16WdcpERBe1h3U+QzI
HbjnC6b4IZg5B5GOj/jbrVoChD8biMDL20jPtG73L9D/dT26W4AQ91GJx3JaS9VQ
T/0g4dwr4zQSlOrRZefZd6Faz5X+UqNolupl0X5zl2rCVWbF1xtGWUEN2ciJXsAr
Pst5OqRKp+HP+psc0oV2cO4rCODkKpxozNxszG20M8lSl0iW/qn/CMwEO1QcBP6V
/LfHr/OCvbwu5VSpqShpTdirFmA+vNNtDobs2UBH03o+sRLUPsbIIqGRwC/x2VSI
y1p1pnXXpeh2AkIKuT98CRkPwpBYMCB12H3v03o+WyETfhY1ZtQIX30NmjSGB6YH
k+J2gXci1g9a4+BrGbR/7PnP4C/Cvvrk0dQggYaCrziSqADYn0vdfGw5Stn94IZX
Cpk3plaCbeQeg6jI+RQByrnjWGtVfvziQU9If3CtlNy5knbfHvvcewYi2IgeoIG+
jr1WPzENRIybrHmuOnkqLNYJk4ObYTx/9XvrPsQe0bfnzmOZ5TnnawPT0TZsXt/M
rkZnC9zqvCkoGrnH63qusOGBoOQbAOn3Ds3IH/zSp2RXpsLLmncKtUrANRsgSkZ5
AbcxPanvCSnytAWmc4BJkk8KGnuoU/HCz4qFnZ1EDiPkA5LUo69wluA+e7AUju6N
41sTyEimGpLrcRb/PqgwrXbnbonBjqLcZDB2WdeA3sB+m0hsQusfK3Nj0WC1+YD9
bSAjacPox5RhAVPfI3WRU1eltmIpmK6hwoOJ8Z4ndccefDvg4dcqlZ5bPfFdcUnp
TXk0z3ziwMACXEW307d/9sWe0GM/jLf6dCMoZu2orZEtazoeac4qVkA/Raj89wU3
4Ew9DPBWzjAc+YEhH7xvKg5nVjIlaXxIcNn1UTK4WPjpyNE6ZYLRMFeaMnT+Lb+c
NuOTlvGEpLIZVhPo0qSizaeIbohEQat0lHSRdmbHoJy1NZNGEGKG2mIbrZJ4pMrQ
URbAyvBocu6VxCYquufpSh2G4WPd2e9GFOH2bGlOqbhn0VYASgmbgFVAtMC26mUO
RbzFUr5qMD8oXsbRqII31oJd9RtKGd5HNsv6EVteFcBjd3aIvZlVzircX7tEnY3s
+y4IYD/0SNMtNUYU6Gg3awET3CcrxvT4rx7BKpr9T6qy/ucZY4WLccwkWTw/8OuH
VU0PvkB72PhURHSP9R1JjSdIwsWoPa3QxTpjxTPWkcYUfh5IRddtJwdYTVTuZ3uH
2kf1sVogciHhazeLsHEHNwx1gdmiAANbXXs2SCGVQYZn0frcHj/6KxDx8x7+9xUJ
28Lnvao1G3Ztw7xSwTPls7E1jre4GpjDo6nWtYJcgjXhJxLJMXoDyn1ldMGqRatH
wExCmQ+BmiJYjjEbDOWeEhHQoP48RUy+8FwovDKRQ6GB7hU74eWbtxgG80L6zvL8
3pZsFS7OgFhXkTTAmiSH6OCs3wMC0VN/pJIIdHz1MBbWSxPASM2iwK1uAm03CGk9
pf0j1WnJBUo7mM6Pja8VOK/T45OQYZ2yX/R01teFtKftyO1PLksrVnEAFTsx4pmT
ghN910tMXeLxxiN4OLc4PGema00TiNRNOqN3HNZHe8E91mZFruczl7Tw7x4tYEzX
wwRAEwNlhc+gmihTzJf2Gtx+8BeujSov4kM5c0Toeki/oDtpQlhvUbcx9J7y67kB
9lu02SaKbGs762b3ZJIF8BpHb3QwS70MZMvMpfuf1DWD7P8OVEHSoM2U1ntxL8/G
W+E99yjJD/D45Ea7E2E8Ak+lGcUD4Z7aEEGSH9OPQvmUDxF+cm5gaKHLkWNQRDpK
zSF9TH98gOV4Xk+iYRlF/+dO/aTdZ2KS3Hrr55QXDIwnm8x5C6+jmaXb41EWQOVK
r4HEh8Cg2GiOzWR/3Ho58sda6gaJXMlhljHePDEi0zpJ9jD3cpZwln2hqY2nRYcV
cOc5mhDQeP9IX/hn5g2Ffs46IQrR4JMHhUXvf4/eFvMUi108+oPcfyotXBaPHHje
eTj72E2mudKx1pjiqiAx/W3/C3kkozABXY01cpAqE1AT61GqoFp3XHBQK4VWkrPM
VZO+BmZ5INeOEnLs3a5zX5rayti7SvuXVPWcrTCinia4JZpfN/lhSIdX+qZGpk+S
Fu1bZjQOY9zq2bJAyMmksbRIOOkdD6aZqiiFnURgbj56vbxMA4b/LfFEydO6R7Bj
sx09W8DdyE/oOYA6uptx73K2UyhKkEmQtId7roXg5S2+suDM9hVYnldORkLokArx
LKnunip0dwZEN+sOCd/HQpbKP6lyzFds1tA855RV0H6CZJsTDP7ErGB7hCR7cMo1
i/0mAujk4NHvLoZQ7R+QyW6+kiJq+kq4iK2autF8tG7rjWm4A7yTyNGP32/Z6QBL
LYQYo5n6WbPaMB0qtxu5YBNPkaSoWPrE7sHU+KRpMUL37a4MSikBz76yyu8zai9u
Yz9mhGDcxHGz9w+IHls0K1AZ2abAMeRnMMAdW0+/eUVgX/OnU3kGTeBJ5TZyG2Hm
1Reey9E1iomPhCcS7riLCYMUv5A6iZuan1u1WWUvEp5y7nfl2r6gsWl5iZwsQefS
mQRD/SdUzpV05luXCNRXGBf7KFjkepkWTw5E/9MX6iM5JKTMfgiREt1iARYImbNe
ApyAOMNSOmCgO7AQRJArz0AdVWO8xOQhe6XTyzT3yM/9lWHtdAfWslGVs+5NoWxo
wPEgj4yxDbIkL+GVUkHzO9MX0vqoaFdym47y9oKbGa8xmo6ccX8eK9rhsaL3hTDd
jnL/r/D31+coLAvgUh22t/HmczBaBWmQg2ilYebhjMuN5IOm1yctHEV62ImL685r
1nxsbWJDKEmcUFWTLKpzYoiGDKGfyrVOmOAvf00vjXWilRy+eVdOVKohuYjzDUSB
36YfkLBI8NLj3Yw5expvxrJ8ZPD8uMq0t81sbX/zyYwJm7mMwtlgVrvn5jT+lPbS
pXYkt7oPQvK0MJXh/Gxc2cUw5u+pN/Wyh34IiklMnXNr1qfkhsyDBNok4XNf9NdA
JokSnAvaaDtVQx0QiRg8jbxqHPMKIMS4II9bd7l5yVpb1+yMm3lePcvn7dFZstE0
G72k8Cg6KEJwyN3S/mD6GkAnsVUrXb7K7ku5ZoYK+4jfX6v4ugMRS3Lpx/3zsTt8
XXWU9481Bd2cOabDMbDEUnhPo8eSdbWW/l3i8DG56QuOxN6ZPDXGp+Ky/Wy9Txsk
w7sd++YidoGpJPMIlx+LMq1dpgFIBnDIHKNmPZAgGqagaJ0tKdU9CzrTKVweLRgK
cgIyQSQGxKOpaseWhmZfQ8MGi1GhWVBXvPyYkMfohNAxkfBJe2EFJbYE8L8IQVGr
6FUrQ4eFqW1M+dYF8/jny232sLimY9OVNZdYPjVANdL6clIVUbdqEQ2aTF54KCGg
Tmq0QTinvV8Qq8rkdIDsPbPXZ2eAFHfo7TV3VZKIIc1dwYXyJvtlq83Dj5sGgDvl
kLDi25tP8m2edSYBZTcFDeeVXKHi57uP2DGFRQU98KCpTfmoqi77cJTkvWYmvK2R
xxSWy400NbvCWwafmPdW3Pisdbd2HmF1hoQwqe4UiUz33Kcl+SNXPrKEzZnlfLXV
Cr/eSmfvtqIDX/0hSwDMy0YrU0QJ7i19fH7i2JXlt/MJNWqQmQLMJ6+ix1LCHtHH
w7Xvg1Lo0MFEAs4QyeBpy7BCfTE+SR2tyT4VoS1U6aoRauWwti1PV30h52qe71EO
1ZV0rvnGUn3KZX4NDWI29M96FtbBiDQtZl6J1yAlrZp/5evcDdsaHqaFf8QB25z/
VJssrT9wTG/6To2WmLJ6OVwQPzZf5NvGJaV+eCfWbVyOok8+vkDRj6YTvVXp7jXD
iFoDsa6DBPfHqovIjMf2vjgeAkCBJFUI4VVbAkDRBh0r9C//+x6HHueBU5Zr5iWe
Dw15oP3G2+QBmhxkvundJjsJMjk98tw6AnNIt4K4hrMY+VxN35GS57tXKkaL/Hj8
fVslNIO1O5+nZYde+dXpOz+Rob2fUMObZncx375dtGte/gttlRi3nvS7EzgdE11Q
FsvguySSTYhczyyyYeMz6vu/Pbm3TydXWD0wj35W9dM/gVg21A68B8VC2qG6f/gw
ayRWgxE9nGXrm+sBsAEcvMGA80XgfQ7rylMsZNxpEccgHpNrC76Byt96Lh/mVtY5
OGGCAjNO/FcBQ3HO+T++ENV/6ofehOuUMc+K0x6/ObosfuSWtGlDmS6Pr/KIWR5n
6bk1ZLvX4PnLpKd/27bBNki8ca3qk9ort8d1Yfkh2u2+aBjAvmLlypM9LoSNIAWM
ZWTWcAUD+CyZueXbQerAT/sxgsDhwuvVJLqEHgCKWZrIAOkIouNb3jcI2Mh1AGKf
Ruh1xgwCcRyJo9PA2027gZ6jxI1hDQ2EKwcZ01voI1X/trWE3XMQyey1UBLPHO7b
vj1PtC6/+PM9DY8sBhhIGuFAv97HhK9sHF4Xxuxvb7Hc3xFHncVgAldOW/JRd7Dd
jhdwBNt/mDfsvDU9qZrlbZERHzeqv27wzAvWNe1k8vVhiTUNYisXzUNLqJqcUWb5
a7MxmOHEviQ7IPvNvVoLQTUD8fFOo2aWSLd89Ip4C6ZzTL9IMPb70nJxhFu6/vsr
oeXuiClWfxbNfi4ukxHCOErKllm84UIVHTEHCkUY6u/c2ZVqetQ6IA8Ur7ACYd1y
hUKp+5o+vVWRf8veXJO4iu4gqWBeJO1TbOLfAIHjhU+0MNVgPmN4Ac3cTxBgOVzI
DGFqvozBqqKXk41HlyDcmy20lOGud1w9sfbAr6zOXvciVXeDHbiptl3ZKB61pNux
R9/werzm4juQ4TS1bGR5wKtAFEHn+6N5TPUDhAsFdIeZjcnU+c1Lgbtk9sng8YvX
DekcmlcbreCpGN6LVVYc2y8oKUN/Lv2tcQhP9arQvIt/yxJYu/xnP11gs/uOn+yP
QN/9zmNmyLhmTOYejfaIfPCMxIROFsda8KwQPUKcoDnOyeUqIdfZVr0GrnV03Y8Y
A4uPD1oCV8AwwjlR2UyQEt31oONAAtZr8/FyvmHIrJlzrqarwdYMbL0bBV9Uo72p
/L3CnC/7p6PejS5RlGHM9mpLfv0wRNHEW8oBUuGPA60TvxTB+bdD9oa4eQlWAMSO
zpmM0xxhKKYY155Pffq/nQ+eBCwbWwJX3Le0MsDCFYcUQfDnaL5LiTucSw6Oqb65
scIhPcMiizfi4y5qG76k/wYtcGKlDgC5LCfhkOvaqV6/gsop51v+z+IwCtMsJjB1
0Vm7EC2T5eGXP6Jc0vsCr987G2C9kUdMdAYLWz8iSlPSN0Y+paZG7Yf15x5jbArN
JKXllsmnbd8uRMR04T/2P/V/UxsjDT8OUdNL2SYfGuftUPJnGzsJyi9uTFCV6yxo
dwNGMXnYPe6zWhMqgo7aph4y0GNkmsE72CcNOAYbL5/a4fGhjbw+cJrJ6HAOtKkj
0A2cBKXVfrLkWuw4Btghx5ChAOrEslP1AtdRs72o1/aBgVAs7eaba23qJCKVSjkD
kn2LvNuBMsg0LOE1mzikYUU/yRdJqka3rRarNYZL4JVjZNcjLsOE+HvBJFBacvii
QavsL08MLHA9azrwk+B1tuWK7pkOSZ3VUl7KgIvSJehgUCJ/witH9pEJlbaerJKW
cDrbW0kZkh+iLK/UTpeaDu5p2QKuxUEbdH0Pfk3iZBdCY3AoYRJigN6tAwePpNJ6
A/SOE8m5WsEAJ9oQDS9H2lyDbTNTdy07dniJc9Bd5hmeyeRy4RIUGuef5iC2hfeJ
1EYpJExUL8dY2FqMxxZJl+EH1gegrSUFQdHGlq862Rw26MGhN9AWauV+TEmiHlJ+
EZ/cVTmh0Ze+kXrp+FC5mja+NOfp/9byL2ckq4C1lpUh4tdvFWlB6wizabVyZsrd
aha56CoWFm+mQbAhEZc4YpFS+nrfgAC11YInTfH+bx7X+66H7w2cOh6z7fJ6eMEh
ugUI8ZT+0LIHbKeJwie/TFoUp0z0EVBj8lMrjraOtdlFQMJoZMCQ7Z8b3d+NSoJo
BICdIJPgXkJ8CvGQf4tgBBLiJgo7aSF+FDmVwxXyiIsrQqS297eyZnjPnw+YonPm
YwptRhFJkzJ1ZXHcMjQllB8M5AskeFsbxT3HeAHLZCdHaA0LqNzY+ZVVRw+5vCMF
6O5+3gCAP8BtkxSntgORMxjgVvKD0lxhCJQaI9nNgKKLqgusnGv3roOPZBC6Er2K
6a2bI11SKudy1UCHvWsDtnopA5YSpiG0Vm4gE2dQPCjQK/SfCbm9yoQQXgwy23Dt
meA96hRzpT4O6Fqsx12C0OIJbci6zfcnEYUF96HfhoXAK8kAbUa/AuhWlhpBBImW
cZdMB0ekne4qmJFgRP2sGhhLc0lGBLlPeZm/bQiOt/7/UtG0XANpJod2bny9uVk5
ThDFgQ+WSlmhIY2W4lKuDvbFWOnmUeJz+UutCHame4h95DzeUMg0ikQ+P97GgECP
U7dBMSxlWvO2miGZVPOtvok/V76o2dhL8wQYc+dWN3oDJcFxNKYlgZxSe4ncOTlz
eGhcHkFvVMWxqcpNu6ebTbRQoCpd15djPhfLoJk9RivQavAClbFAib4vD8/htFeW
SZFRDv0e56rTrykcpdx7rCltPFicAdgytUXiLjHiXPI0oTM1Ty08KZmCpe0igG85
man2J6mw3u7OeFSmZuLSmB9QwmlVbhNUB9hUrNgtRxNqxaFeYKWEd9uVzUmBRnI8
q47OiYb0O1PxiBe2aKpxchggnR3CN+gZH1zu3yU/zn44OPPvswd/7uyyOvCQZZM6
fswgK1HfvvWzH77GD4Bk21E36fO3pQb9A4ckufkmwfcOr4Au0AB3ty16zd4ySK+w
ojbxVKp5j7kgd5PZ67m5pdEYeFdquw5eezaTsNmsyrGlgIHW50fW0yYhRpn4w7Cp
VU8FqmKbwmULT3aByLHTlbtVjaa4DG0/PRdTQt39EJzUQjq+K8fF1r9sS2wbtqdF
FAa/jToU51q3XI9IVHsMIU82JnHg9Op6TYp/WO3sxn9H3urN26XLg+tUlktW7X2j
5brXbWI0cnbP1Rj19Z7R1jbjmeO+WHlCXoZBuG8Cj2f0SaGsN4/WH/OxhJnQI18f
tOXSxSPzD4E7Vr+HUg6EIFgxWniMuYPLvB+1qmDR6c3AsydQ3H8LDX1oYF8xPCcJ
MBnjY3oEkO3pQcTyjz75NsejN9tvz6tbhKENvmVe7XaL2mSoluol7LLIuCwmjHfO
Es89tBCtwATgLk0Lh3cVe43fotpRHSw0xX3NHb2k8VWv+9zH/pitWBPhf076dFQr
2bEG2H8k5Fns6KTQa4nhfUSrO3fXYszfkTPNH1n4bfUnpbDFmak/rNikdiDvcXDf
WbRFX6BBON6DQJTO16ALRnLHFidqyBsnxyOnM0eVFd8YHiMY34ejYQmmUYO8K6FK
eOvXZ8v9M6NS/Wfgk3eFPZz9eidrWxfO+LePG0+jL1Y04LiQWzyw3ztsYJ+U+IdW
86HWYcdgN8WZP9hh1oAH7C29TLHLileVTYdNSwqZAXhq2cVTK8tvzGgkmv+gWjM6
6Ynh3JctsTGQfkhlTK3xFm+HJXSvpvwoPCzhq3OEnKLJ2UV4G4oEnjyLF8/07O3s
MJLiKyyUzCFKCEcVyIN3hCls2LJF4TKzbeM5micE7Y4Erw4yosYdFpz70Gw00z3K
+H1zjJfTijFuEozgzY+9ovpmF8pLwjtLP6pP7r2rOE6VDEBHxKDTIIKy0jJWHBHv
Erjxybcd9oiuzDMQVKLsU1Mw7hni2YKP96CNIRv57BakkTNP+zhAZjnWnU126IQ3
63HyvHr+lbVUNb9wFGZJtKfgN11z0kGGc88mftgmYp1Xt1Tl3OCBnyWXf3wBSt2+
w2tAgV36RUYg2SxbrZRxTQ9JNJ2ouZRYjmUEzUJ85GDCErdTqkTwuja+1Ns3aj1o
lAd+iYu5hzNMCXQPgIHJJmAK4mH53nuc0/Yxy97GIXuQ2Mx7Mz31zy9A9ZBSgr+I
xNBDkjFD5Aryvp3XZC/qxAQeH0Ebc7P29PvRPjXc5reKGM0+tiXy3QXsO1eu//r3
YeJhC6O87oPD3PfFXQPqgwFAIk2dYPdRwVr9DXS9LhDvuy3RxpuPTAsXzMrR+7lR
adxkDtwBuLGeUA0G41BSEWQ7t2Qr4BWeUh8lfqrnY7kzn3Sr0PbUNoQsLWhYrFus
VpMT4X6FoBqex8sK4EZMNBb6PZh2Q4kFRuAPkKpOGBVouA8mCnmj9l2BSwOohpDs
t7C7bbkobHsswgr3rV7XBVxmAyC6gcQtUis96Vcp6M7eStfkmETE4AwcXI7LZW9T
Sp8ua5JnXx6tz3HlbL94pm4JnDTwTtZoMUbebvlu+MKftm6vtHyF1APPZ844n/4t
Jy5yf6EPsbgooK7gm+IjJQIIKxwoyz6DCRHADUMhjFh5xuHT10KTuvFxQ+CUbIt8
NitTVU64R7JTTh8uJJ3jgjJJHwWo4U+xP8ROhq3YcfHrWsIxcYw5lCnjScr2MzO/
Y4l626hqSfKRez/gwLcOnbQ98QBOJBZUoZFR1n1DSNsT1RdyJiu77Ub4zNLBsH8D
G0/SL8/7fRtwQeLUrSUfJTBVIKBBUd+U4eQAqLMBIBVU9LRDrjsJlhYA/cAJQLCJ
LSWJLrNqfqjGn2lFVkh0gyOSif3aNhJQ9d+ayVNX/41Va/EGUwzaTzXIDb6uAcSI
65xIzyzy8P1lE1f25rbOuItXcFNK3Jg5B0yRbnZQEFPPlc5Trj/w38yRpP5WTJwY
l12ERphKTO9ssOioW9wwFVIYViJCJXc8HyHpO1nBxZit/wckxFIYj0a0+eJQqgvb
asn6cD1IPd8+e5YYqkINBhqOTmaJBrK3z7CURBVCnpuk/4BeHRpLJZhxAgy+WwtF
ccPJmL06AeyxOCwNxXFQQiGaUINqYmwDL7h7H6gnl2NRCgQoNpDeWv4FKFxBIrYg
E9hdZgYrLvRClVrPAs4/v1p8Z5BFE0+DoHzlk+KkwEzh3vFW6mrW2BzI4w6zQF6g
ySy6aW0jjitpjAgiySSPqV77/GHYkNlPxhCJzs5rivpUr1rQpf956cD22bR8VYsR
FmQcexAZLvdfIPS07eGFdb0P322oFMPpnccdH2erT+ZvNcjVvC72BoFP6+ICb3RX
EwUUb+44xmXbd2pMkD4WiTnhIoabpTO1Izg9yzBrde0WHqV9d0E688cjXIopfvnY
Z8UB+/6IMzk40wRwyI+43ciaYg989/LRqc2jRkAkdaB3N18Bp1RNk1ohzLlJ3f9k
Wm4COjFM6JpcKaJy/ZV0IT0AQyXp5tTSOfyVDa/E3BIfe7l5eG6jDRPIr4U7PviO
1Kg5M+BmfvxPz71CaAMo48KWE42cTMk8GDRUmq1b36X+abiQYTVNOMG97aJ/1OYa
r9FGW9Kz4fvMMLFdsMu8kQM0hVHPL6O0TnsmnPz/3ICpNhtqnSaxZsl44Fh/Z/C5
GXrisInOkNkTtYccmx2r0nvvAXjiAOl7IU3s3f5zDPV0//qNdEXd1llIcLr6Bfq6
JTfGTs8tgVU0gC8ih/X4fToPVegocHk7mqo1y8M6IUQF384nbd2AEC4GoihSAFRj
gwTzDw/X6y4FBJF7d2iKCoriG8ucz4LxOKa96Az//a6n4+wP7cUpF3gYc+9ADpaz
4yG9bjasrjvGxjyjdlARoW0Qn74V5q8sMKj9WznvSiZ1u7ccQOdqE4+9lwbENVpI
4WBcjbFoZDyq7+PwS6PZOndg1poAnhUGe/GzfOlr1j5rgIFMEaXfokMVvF0J3Six
T7K/4nqi1jcYmhKfLYKB41YZCBeirE9V1LFja5ODxtm+a36O0XRC/GwuIXfPBbQN
q+CeknvJh7SWx+46G4GAmyCyo7vavHxoBJphyKZT5P7Bo50dW8uop5e0Szk8/Nsm
Jh2yH/3OK3Oslqha9a5Lz9MiA/2rwM54H0l03vidJgvYj2dog2Y4clYsqms7zyN6
Vz9UMvvTbl9CBOGl4R3A1IFwWWy4ag36+rmgUdmwtTd092PMD5hp/v9PiCYdTI0D
5XXbhdu/e7PkaPextW9znD9vReRmsFvSdJ06ykfQk1iPpi0VbfjZT8j/CJGiah79
TY8Riqdcw7x4wIZ21tO3O6JWOPgwYe9MG7fYBikbdI2d9sxkhDXMMfnqd01dAc9Y
vB44fDIjII6ESBvB7uBi1LJnRU7QI6wSTbeAsS6JJLHJrP/7iebDfbrgKdmcFzz1
pLKqBBEilaTdt0HEAbTvivY4uuG+KLWawj//d0fUf5UPfCYVlLHkgjO/LNUYt8ff
MqtRuYOTpuuV6EpJCqVp6XWkz0IjD3YoYfRdG4S74MkFe1gmIRQVqKoDGyrMEocb
u+zN5fz7gv8QMK1ot+IbnI5w5w1ofolnGVyN19121GQVPkhhMxKZAbZF589o7cTR
k+8RbNgTgJvAOF9E8RvRgf5qUOYTT8XBY8ftB3qKBOZrbeMVsUCopLh5Fq+bfVa8
xvAiVGACa01IoVWeeyY04itI3ocfiyDcKqD5jTOZP5N9TfI23ziTdcQqMBrjXz3I
6AkuWaVZkrDutfB7RnW9qJ3z7vJ3UdjfjSigZd7XuS9yYpqvRfmBTUCW+Jasw0te
YN6We9M1sdDX1z/7RQjYScHsbpvSUElq3QThKDu7uc/aIQ6uQmeYNSE1xltSF1y7
gHocGPyMfGX2avuD7MZet8e90sTbofNVQJkBKFQQWfu/rXdAQRQ3T9R9SlZq73f+
ZmtD1l61W8d6gfquRxsfGDDkJZ8Z0QpP/1tEwrWNdmjyUfCUdXHKA256cnClHFAn
zUDi46587MmVR1RBwLC0yaUkjq0mbSvqhmtkRJB+H5LRADQhmgkLhpz2XsNX3JsH
huL+ytvo5YMcEBtXOKYkF77EDEPdEUql3WEaGnKowkU5iqLPX2gfKzardxR9Xuio
GMP0EM9ifJe3A0mPTNJOSQ16OE7zLwhTkrWoNLGP+2Qown/hJVpigKeVSyKeS1+F
5It7ZmhxgKb5saJ0Oo/OIgBpdBdLM3BiAYtnBz3P4Jb0Py+Kld+/o0jP3x22noKc
2pizbsc1l8K4f2T8PDGGxffvB8kd4NNpuPiYzY0QZ9+l0+DbW5Fdm18zEG0Tw+DX
pB3nT75XEG4QbZtSenctxPhoBxvv1SfwNwrPHTxcjvsRT71p6883aRKRjBFBJ8bI
OI7qeZsghxYMmiRMMOJZpFmvTzHRvCmm3ywAy4FJ/9i5G9hSRYvMGE9glY4CxJGJ
fxqAGqD6/cKY5DBQWQorUn2/p5YhnLTofRnPlGtojrGOkaXYFl1yz325nExfgwCI
GHAgaVH0R5QKR5xWZRYODWed0oMti74WBuoWc7YNyauVYYnmBPRrS1Z2rx2l5tHo
sDIZ4iGmKLbRa96zBUMSJ2mfo94GXydyOptq0JkWfhxiFLl9QmppNC2NjGfp+7cd
G1JHzZUWjH03+5vohuENAB9RnrkwxfNhtivcrO4TfxdVAfjwxarYq6Hs9IeZy0W+
gVXgD/zQ2JgfBPylzb+78gSPcus+LbUZvozl/jsguH/B+JMiXv6ATjiv0h78Cn19
3a2KsY5lWlZK0vHH4mw3pn7VuENZ/EyS+NRoa4oc7zo//VB+HxPttk5Bnc3oHkr1
tIeIuIYsCPE6XY+0GomNEH8RrbgbaQSJ/JBhIu0zlfZune83TgCvO/5VRu2C1c/I
YlXhtOYoyZgdMO+JwLwMrW+lIWs01pOlXRknc71DzYa7nv1cg0YtgSYkD/s7gb7J
2MLehRqRpEK7AVlHE+XWDrNX8jNpJoY4yl0TVdlroPXZq7otUCOPW1cDYSQen7DC
bARhmDuyL5teXTGG2NQCNRBAsqIap0HrfEqzSUXh0lrmnEf71VYF7X1EkdXh+gsD
O2Y6jWB3sKaO4wEIVsrYwHuX/GxC5Nyk9OZCCS7ZPt7G2mw3HD1F4YbNaobxTWTH
J+NfmbHDw/DmRDxVVJlGvbaaErZbICBI+OQ0hOcMTheqXIKwdZhSCwrDxP9llS1j
SqTK61QBr4rV/CJcsjBTYENQ+6uZNsINg/0InXvGsx7oA2NVAaWQCsKMiPtlDDJu
e7ulVdRkK6FbkPWWq014KbHLjNPyv3BQ5m8kmgbDI6PsNJ/aAzhodNEv1EyVCCWd
vcQf3jhf98ICbzKBqmEOFsihjwShYtMijZV+SoBPvzwH8/6U3AeHaDWR0lJYHDPn
lkk52SFz/FjY9e+8fnGANphR/1FLkGnnMfRkpH/e1jQjabUklhEdDIMugJdYSRx+
qpc5PIBWqCcMrWl5vQaxyCo7fc9Y5Cizl+yIgo0ITbVb46lGKq7LMiD7koFZuzAg
Vdt7zX+TYL4+MQ5ZEJJvGH9Rj/k2pSUAgUS+XqebxEFU9M4nkcC+lqbyNROixRFA
D2ZPRQZ3NqhAGc4nZiVQ8v4DVHZHBv4el80Boq8jido755hMd6NdU7n/zn88bPKK
PV01nmyl+UjcpIw3opXVlLMtnB/X4bzNn7gy8rMxAD7F7rAXj8ykhZk8egW60Yk4
OBUAaOvEdaZMXOU3FVo3SOv0URFHv+hmu8w1w8kz9FlanmLnzOklNYZ/koH773AL
gnwAZFIRxE5zrDRjUABmP60M6XRXoeh2XGoa2J1wAfhDC+jswRzl8AUInGqoABOC
DZmqibeVTKfqoza5vnSoaatR7m/J9pLXtpp8HV65lBdgogHD96O9OtJTkE7NQjeZ
Tl/hYZ6XMnuz/bmomnhiq1qkfNyH3YSs0j4ZlLs2X3BrOpe6p7Gebf/1AXX7BIQQ
hELQaiuae33LHmzibUnjG+0zFcr9esxV9kzpoU/YFSA4zZ6LeoPbos6vfOOyphzG
8q23/yP3Xss08w/XkDvq8aClhNHhbtbl/zznUhKpxQsvPfXoM15yVyoW2hRRXFIi
0ab32uS4yHOn1GwE9DZfpRtzDS4fQGRVkUOyIgOmFGU2n7NNk/JnrtlyBwnJOsfc
lzgnwbg1HFHCHytJVR9PzDS1ZP8C9henG9qBA3QCM6UuA5X/BwW0NfMa0cSFjc4j
a4Jrv1lkG9gsiiBSLSDo75g5nmqtCG0rEBubBTX9zIzZ0hmwnmJf1fNIPhcW/PFt
G7M6tjyUVp2Nw6lt2aZdD3tu91Lo/FPSoLAwUt9Jl9C3kJjsxqs99DSSnWFkhZQP
JigC0r3tUecR6v054X5y9UwKbFyWdkzXMErlLLvp4Mb2LcTzRJcmpyZBE2vFscex
1Yd+eDGnOQOp3kiDK2s0IWqjdCo3TGz1+rWtHoZuVvT9VCyRR/XoUY0PcMD9URDN
tuHpUc+ypLCfMk7fkLjGgJLnfCrGWFJ3qUVCikMXPYGa2611sbwzuDg6owO9wFp1
RtYlfW7EiTYua75tTRxcqM880QR3Poso6z1Xf81FGSid1udbO7U9I679TRHxPYJY
rW2tpmoGn/CgcRdDSksOTLHcPv2jXWtv0Bb03ghNvD0H9vC3YpdWh/rriom+AiAp
bsyl9TBqoCxJ67oxOfT9abzWNnn5xURCEWpXvG8XB4VJw6ZK3jQ3W6PtglEn1E9i
FEc3z0Sq2XnS/2Fq1AQvwCFQiWVbc9ik3nDmeqKkYGIZ1B7QGp6BgQyR9QRqqsuC
vD7peU0Rh8MYs9kBU61evODwwMOvQNeFLQUii2sej4nXhX7cFkqNQgT0FOntq0NC
dQMGtCkwUW49UjmZvyegKbbngpDyD96MAsszNr6Mu3/ANFEf/wVDSpKDbntjBaC2
EAo+axEd6leDx0X71ntpYgc47S3JyaXnguA4z1oVjS5akAtQqTcH19EJ1XnOysm5
+BDD3dIXtcMqiCHIY5dae9aYiudkizdeQeWGfACsjHCS+U38MtyFp7lV+Cbi7i/m
J50hXpE+CfZ+JJ63cHv/tQt4+eqjyXUzV/VbsGqtKWdNqFNxz6oIf1hHAeY5l8YR
/JuBBfpyiTDysmWvIJXlQtBSDw+xM3ZdiQSBPxwMAg3HFBRPX3TJ1f0LElyrx+Ts
7FZg1qwJyvx5FpVxW6BizDawAaY/TmHIUpNE39cW0M4sjSazAB79/Swm8XPneOnG
Ipxyxz6n3AMbYb28ohXBnBpoqiVlKDmMU3ylc/BKIliZASwx32X1AQpSafIh3RIj
aibvPLJ3WCQ3f+1x4jqH1CZTH6LSi2FydTjENgw2reiduR8wacUi6OcGMU6s8DUY
UF+ynMbQkCdYBqe7iz/pBgyb6cQaYQu+pfSAXD1wBMKvYNK40cfGeXsHpmmjS0CT
8SCcPDcQ2r7eFiVZBBLWyVgSp0xlNir4UJ87hLWU5tlqEz1jF+SQEAJQOJVXV5nL
t1PpZyFOvxNHeeNvXiXYrlzRDTDbmkKarBwwboGka9qaFjRr8oMAVvpnMe9pG4F9
+ZpGuA19iAr+NF/f4f2+OnFwBKpEzY65hlGTQTpvfYrT3pEKOAAX4gCga7q0CfSY
KiGzOd9t14qsBoVfml75CxilRLrsJwBVJm3e2G5whvky7xNWwTV8raFexTCVqIbl
1NornYfQmEtWIX3Zck+i76l8kE+JdWwoEPsK0gvjTfwiHRXdsg6TP9GADSDYKzbL
Kx5sHb5LgTsZ8qgi7c/1dizM+RKrKLcaGOj04iYYLHQy8sbmjpTMRqAxDnLQx5s+
WmZRMhD52IUwC6+OB9sJE5Wsxi4a8Rgv082oBXASkEvYXnduJ6j1iGnU/T0ypanG
Rb8H/jdm6ZNpt6DbF2FgRGBbfFTxNVMSQe8apeJ7MMQWswVILuAGj/yywn57Fk8k
ViyjdAMFJvwf6m9Gfss1yGD0uA/nhgZOQbvL1O9SOj1V0f1tOAF4T5aSGnMBHTE0
MXpH+aSaJC1VcECmbqMe5Jkb2qIOiVECy3uL3dgDfyqboR+tN08HvQm6HwSFy5Zl
hPxUvILXsJoXYBNooCcnZ8jt4c2RuWiZMRi0TEfSoypBcEVBbnbtyXm2k6OiqLXS
c+NbWUHDObPrnS5sy9h2knaPd+mFtF9fICvGMB8Up63l8GdBNYxA4HXLsKHgsFqK
rMUlQ/l3yDUe/RhicyS2FYCo+qpynv++nyc+GdMzqNKPHbVgoDqNqHocwqx/8rjy
eVHbQCIGEqGdKw+MHkadyk+7PNL3Dpv3pkMbP7IeW5F5KfnrBCMQsBa0P/BIg0h/
5sPShP6BbqU7yGhV1whJWrr4AkkW8C+3x2owBIjpVoXE89NkVH3fX2kWrX55w4NR
AujORUhDUOOQAh1A0Cmqlm9bzFeww6mznvVkyHAYGo+fQqbDTU/hq4wKvb8Jh0X5
eoTVc61fZsEIYODiSfY6NFNzV9breKklYz3i/gaPHmpmzAGL70Z/cdfwXwSUegrU
wl3GNop+n+g8SU5NYCSMidyrVcmuI9rH87eFPXm67KjZUeNP7qG0mz2sdi2hS56l
VRnjnbQ/Cn25H8eQxsYUXs45Gyfs+wrv7tZf0GNm7LPprVRpWSPZhEXgvaoROfnS
eE9T90/DtW7OPhcYfo8So3hBXY7WCCu27b3EthzG/yAY2pZ/LLa+ZnJ1tSMA2QUc
bg7iv6qnZm5/X1lDSBlCCH4ChhhrTacG0fSwSGYQ/5qkQXDwnnZoqPhAP/c1KZwm
vHHsvbgjeDiNDfuse/Oj7qqp2iJyj+mwrSaBzphJgxv9uVzR3RsceEV5nVCqF90C
di4eDnddzQSaSEiQQYxMKY60g7BbKmcWhZjaN8rf8egZ0M+kFalR4nw8UDhlrO32
jDxEgzgy+2VZ0lMAyYwHjunZ18WQhwVZy+8fqkHHpKD25yjCWdGWeVRp8k6p0veg
mAWssz6Ju5LS4G1m8m/Q9X7MV31LgFXLKB11EjRXKFHBcVFFetVa6AHYNfCNpK1o
yW0VaQuOj+aTl5wZlBzX9uaU9EHCoCGlL1QFKLavGYvGvUDnREaIMqnOABPESh/h
ZiUtgTW+hZB6EfO5sGyZcXv+Vjn0Qe7O3Ty1WvOL6wugL3RimyaFUR8svtmfMfkL
/7YRQF544WV1d1khBRcH5wQ/RfalANez1UtiK7F/uzELrWghOWV98B5vcJNAgg80
Kr1T1kUe/MCNpiO/AmgiYpM6OV70L4nqMUyFRiVqK3kJlfjrL2EeEV8GxNvdPw8x
bjmi8QInE5Iv5SNpdiJbddqjdFGVKTuDwO0yHA713tKM4xCzYnfoW30X/dwfaK8A
Pow8mWn9TZRE/NSr8kW5BTIBas+mI54AJKgT3HH0RWrN3TTjcPnOkMDrRsU/2Em5
Ll/bQYHcsQ3l8BVpDu9m7BVIQP8wvHAhjtheMGuuU5SpYi3ijU3hPQrD3tp5waoW
Ue6kxOuFuKd0hNtRS3u77sC4I+Bbg4VE3Rcm623b0K635hlpDI0RDcRsmV9+6zaC
VwpOs21+GWMbnriIt50ubrK5/xs4w07FPPNuASeTUeyaoeAcfmSi3cncBXIS0Q5e
0Io233tq+x26hrwtpPn85z8MDEh97ZSdLEhD9rBy8sO6ep9lLLDHCIsmXB3YgVLa
kStY1ch8shlfuwSRYaEVbpPzTSgxtOY4yBqrQjgtjRqEsYvPoMhsMR3Tw2MjPlxf
nTFLBCF+9sx2HgsdSDHKNuw2yGTzXqCKw1iIlKSAY0fewFap8IXV7FHGgHIHgLtO
Yqb6R6DcywtkpPcG5wcfYhfRQETCg3v0v4e/rL4LNcWsv7Uo+D5wgFMakQBsRmb7
8zvxKDbEPkie2t2CjmMpVy0jd0/f8w5hd4vhbkOzEj3W4N426xc+lOy4TSTL4kll
HhsS25Aai0Zgoxu30UFbJrOSe/dbjevQ2oB3oW755z5b7PaupCE5w50kFiqBOMGb
I1oqmIyHjEbP8u1IVBes4jIvwSAf+KGh8mVC+Yo8cXTeMfYKpt9aHQxYjzrt13/J
7A3vLcXjCZR1HxTvioimBr4xXpnx017fM9/Wuo28MlfUVJnno/jzXF4UnvtMy2b8
LwCMvAZxeaBnm0YW5eUOH2U7WDt7crxLZn3SVCoQslGdETH11n1uXTHuALQnjZxX
Doxv3u8H3FVVQ+crdJrAnzPuMGRmHgKD+PiUDs1+B/SpgR3jnhwXUAhRBQgt4t2o
fDuP6rjrOnoyKyEtoRkOQZ23jAyX6acDhkUdNghpjxiSW+tNs9+rsIjNCNxmpIiA
1OqdUwq11n89lfDSZEDBCEmfeIL0SCKEjyaGucVSkO2ZtSb2EksLQ/LOuo9gpWQL
gWCqyEJJ/VjzZ2VSavfvytCL5IhXqJyivFm54i0Y4vbGO6veSps3wuhB4FSCFVnA
tIPg7Sj0WjqfEs13as7wq9B22YQ32Xtu8UR4fl24YP5zrSG6YkM+TvFep2lizqI0
wU8P2jaAGFS3QDfYPPuGOW18nZYlFE3p6t8Ms00/PKEHarS+2wRSSlMGLzAzJkmK
aWuxvFtpuS8TQUC08AQGkRo7Fn6K241IsA5AsnxU/OaJ1PZmCXSnDueYxLCu32It
/Ux+kRprlsp/XpX0UFkK4h0iXXXyZCWQgYdhkcbNr9NKaWz71Rqai6jFiFa6vTZy
cqLyZQCCyZCB6fNRILQCsBBEPpQcrwnNlsmbslVBzhemdZqaooADUw3KtbVGtt+1
10dC83hcQxkXzZ0BCx5HkJDRHg3G7o9VJydJheF7tED6vuVxjE7rzUtOu+Vp5iV2
5g0C7S4O3PMo+MiNrAEMpiPI52mcGcsJJvKDb3wOXs+A8vDXMHUJVWtNNfdplgRU
y6l2GMiuRzlsMVQoyQ91VdIBbrKS1qo7BAr5a/TA+D0bqjsz+YBj1iXmddTykalv
PY2srkf5J4odIVAuyQovRZDpVOKVDMcXXi8RD/m12myE/wpkgrgxvzuqtuYTet0Y
ZWlaXn+otCPuMcBxhFNDi4YyimqZOfjZt4bW3CIqZ1mmBBNnp7Eih0eDFiIGDhm5
8cvRwVPBklyWAcNJZN63P7plJpTAsikid2bJt+HrT1fHZLb9WSVO7tT54pu7hg3v
aMCC1gPNs9kQqFhsZ/sr262g1/2IMj7FzM0Ti0TPCwtyz019M0Maf76mMcisxAcd
hnzbMa6B26ac66KiNGD5VozPTubApBQOqmkvHLesFsQ79NiqnYK+zN83XqIohSC2
pD2vy6cftI2NVnVIuxNLLRg/MxhBg1mKE35cSo7I/B7MCB8HfmKIXR7kcHERoiEm
iWJtEg1QLf9NV/qIK/36Ukt5CbDgDBBEerblShKibILSgqljeDs3NBI3kXpCi4qV
DCQRAcFJkeeyrf9H8pSKJCeLovL1RtYgTe7WDAwtvn7hX0jsKnAF5LcjJ+hAeRhz
ykXPLlK66h3ddVeGADTpdYYckgEX72sh8iHGW27SnFEneOdKpkX3svNtGfM0vzVH
6c8m/Gt4hA0BCjQiMAka2c0U4PtyZrYwbUi8IOAJ1wG/W3Bm2+20Uzzt4nrqKn6E
JPblJMRWyvrgVhOonYbqPdoj/ogp0xNBTi1pyoTra3kLx6XKGhQ92NQac+VCa96Z
ES/PMOyWKnL2Ca5n/ccdYxFyXqFCZ7pZsUgLUYDlYSI48j1VQO5f5Taybibk+8Lj
Ay/4bQZa9f63eTG4/dBgd0JukvE974GV/3ZPV2omhGfn+L/vTAltB0bhN6aePxF1
+gjEIYWWDzwIfyd/1SZ84+rVM6c0oUccYhjGVnruiKN1La3q+5q5qyiO2ipU9HN7
kLVysCpSQEC/fYDsxno4ssMQ3CR1lGqJxv9UEAgrjI93Cz1z77NoRApcUt72YcYY
CvSGTKm2HAoSuGzlrTa0IpSwUek8sW7OQQQbjFF/tp01xhSJ5O1zAtfrHwm8dB9N
yX9I6U5d9RQVzDHdjjyeUtR0GLnXDjbFQQR2lJ4rrsdtBpJt3YkUdF5lpatncMOr
1FTpLful7z/Jt22KHWMhIGwaE7hHFUJR/Hxm5brK2e38sjsxg/J6hhePXYZI5Ikc
7FQfna8qrTO9KtBFWGR3bUgowfPFWPEM8/g2xObQlHC00niG3hEXbq2oxPrE9R9S
Y47IfjqufzVQCqHOszCZ2L2njkD45pRJY26sVdMIQNdjchOvVe/ybofVvQO061/2
4ghdxdAxhMP+1eOdQk0MhvRhg1yOmjlgEjvboYlGP8G63n7z565TAzBN/b7IiYEr
KAF3iox9w5JQZ0eALGzjBVhf2L0eiOnW/hBlfbCBQWRifQeWOhxaf2aa90QG05jw
+y7pGvEPTilT2b5hUQhdi3WBBbNzpcjeSxkJBQYM6MxOz64BMsTrleTNrXOK8BMH
ZZG/+FV4g1yQ2mVVKJPmjV0fG7FgFRwBgQYxcrhsRhTjg2La8oRJJ8CqzS42+m0j
nzIl2Lg5p/Ysv/6kFGSIgvzF+J43/QTpjNYfmFYT5MpMYI81inNq+ePMkxw4y0j0
YMBq6aL0QugbTHe/KSnlKpApUuFUBVoHuk98yIFFqO8Q2i8j+ew6FcG/FzRRMNsO
T9GGWRRwNyhTMJkLc99zNTXOquII1kS22yI3SWdxcYhHwe0/HN05Y43ClCHbt4bL
ExEaaOIB4tTySU+ncjlJl7aPJkY1MtTlUoq6Z9RuCKWm7Wh5vFrFXbPu/ntx7rmm
G47jEP8hzuCfwmgozau9F0Ih3HRliFA212l8B52wGQe2fP4Lv1aJ4QrlB2JR4kJi
E+1SWpLbXSo6GtA+Eqri42BryhH/4JcHyTzZmopxNmUEirft3H1yc2z4AM3uiHpi
Q765cVzjM2aBTxleI2DqHN/4r5BS6VD98yHjNBTT0WFxgFwtT2Iz9+Yc/PVcWI5j
8QYSc9QKJZUKgf66w+WvBOBluHnNBiwrkQeeReL9RN7/jgbrqkPqvOkPg/4r7Kc3
98i43HwVi6/SPnsjZ0EbX8b5ObhNNA31oFo5KkIK/u5fBneIcjU7xQDiiQwEsONr
9bkhJLRZxJ83ZIvSCXH6/J2WiMXFPuMb4IheM365DyI+o/QQqbbbpvjlgX03cy/M
Ajrun56YBpFrV326Ra8doTZlzwp5xlg3Sbx0i7A8fRit0Ri8Ac4/mxmD2k3YRyuM
y/6gTy1UmA5XcPnw7syLj0EKvu1Ye1vd8hwFhWe91VmNWwQED9iqXTDm42AQKdAU
02qG0oGPmyDTRMIdXU8KhZhUmoZCmOrUehA5tGx8KUlf7dUEMN9i2J36EJ+BRwBP
P7/zxAa63bTYMYNaS03nItSfIfQ1nV3vWXI83s1O+u7fPJJqTnpWSlYOldeuGPyU
anZgD2EGlvBDZawgdI/YaPjiyhlLxiZggMjhtnSlO10WCWqvRXzH5/74V7I6lnhg
qgUGfbfpR8X4nW4q6GQFhjpjOpcU3sIoQ+pOyD76wMW8qlKd2sGw1dwEG+UpfnGl
VuDyAV0O1JzOnRIZW2uphvzI7/amqvEUyJEppYSO7LDL5HPnwzSLkr2z+VijJM2s
SRPMhB6luWM5sMZsT0jhjsUqfDVqFjkCDyz4OkueSb+cR5bVScaLqmX1zn53byye
ADKwp+/Q2aG5cWGkp9hSemTt5FrreF7I5P772wjonBODyQlqYTyg+ArH52Ec78Rq
VIhvXnpeomiHiuCSqckzn5Vq6BVQBpJBTliUfSme2oCQcxKipd2UAKaCBZGWOxCp
orrgBPiB/iwIjucJWKaxaOyeuyBLSUp2tlrC2tdUBxH1nIydfZY1e141fnjTUXwG
QEKdsNdwnA/NZsvzaJZQ6nZDbyX3AeHLwj35gSdloofTzDE/0XVqQPeVxhSU88L1
KyGRocmQDXTunkMke7en5wpJQRtodRkVHN7o1rt4Zquc54z7z0Ammh85EkfMxd7e
O+aqSgO4WlB13Yp9dmw6RPGhZVrU4kWANNQXThdbBe2uYlI9VYNDsx8yKa3elKYx
Ss+EVXiYViI+CLYFg7ZPa1Gkh/OV0EXlB4W0840P0HCGkks7wZ5LKL67H1a5KzMQ
1MIWaDCp/pirOq6eFDqnE4HzGasHSOBQXX8aMs5am2NrPtor5fr+a680d2y7rR+L
XPNKXzCeQ+f8qPtw8tVpJZdECMfD+900iKWNQM3RzCVo+Z8abMZ5Aqk+N+F1ww7Y
76UlZT1byd8hElreMlOeT61wcWEzV2GwmL159ENDvTf/aXk+TbSsW7sbiXJP6tJF
HlI2hs1NXoLCWKLkl3pyvdSkSrAxqV6d8edp7YSZm/yx4BbLiZxSDzv2ohI2QICt
C4vxVxQGvNd0GckvZETR/Vg5fS4b1O7VwZtd322feudIUrqibaXoScwtizwbmTOI
/ZFiwQzSu2Fu9GsU/8L7oOeooFj7Jw4UzEI6LFTDdvbmsByHJwWb2I6eSRZABWYk
6WOmehwfGbsssybxBfdwjpSIwJSxn5QgzSKskQZlMW1iykENDOqWC2lgJLG42ojv
Rw2o47lAFr2GeQM9GGMNc7eia9UlC5LKuhLBNheNOhnJGuAuXe5EcpYtTNcwN7Au
AvkszRqqafm7BM6OeZISsi8Z9ghDtiV3xUdQJQudY2Df3/z9dspJWGnBjDJXulnt
UO/LeHccYyPFi8gQi3BTSvaLrm42ulLiM2RTb9QkOR3g/zRhOGaMKTFo1j8lQbX8
epZH2VZpcy0VPj4bDmmAlookAzjxu5SuG6trUXnqOQsfRvJJqA9ANIKAJZeVwKO3
cV5fcT06hnotu9Aa6AC0VAJc6ovPyHMEffC7ASeiWttWMhMvdhpVsDbezyQX303e
lVsgu1FMbndrWXn1lo2dbP+AqKPTCtft/6XL25zDy1tvju1JTWesN4+4w2hHWHu7
YLFXL8C6AGgouER2Fju+7dGfA0y0bx5g/9x/V8yViMBuNK5npqsVQJQgCMwjja36
uZOTYfVGqnIbMc1oIztLZ2F7+lNO6KEalGSdY4STcZhac7R1NJjHzaKd1P/tNqUE
CFblLU9q91tVZ4QqwVbG8r8DokuK3uKuhP8Oys934pXsPhcv9cgcYOahE6T6voLx
ElFJOsJRD+9caOQHrgihldlgN2KX06VcbHHMm+To+/NWELjeN6XNPwGg0x0ayQ1R
5FLYc6LMiGmwx/Ns842Wu2Uel0XQyNNBMs1B0V4KI94Nb4GJVJvaWEGXeKiX+fNO
/vYvOSyuqmSu0eTiNvrUCpZk3kRLpgYBRb4RCMTE+UWqvkA+o8RTnFV1QHAxHukh
t6SSaV6yqsLSpVfsSnypSbOUCA0vBJ7VG46HbT1QpR+tVUrByNbm2k6QCUnDGncb
gxJGUSLPLBmQP+1ekAZ3FQwO7TvHgVlNmxKELZi73q3jkEeb0d07ohun7idxIZ+f
HfGTOnKjGehbZzuQ9Y1+s7JUNZQNZtM0PPdHuJBW1CWOqZs+YSdbp1FqeFKNnwVv
gy6r+Zo/nSVjJHJXVtrYQBYM4XvoUXU7Z3bzF4AEQFXRmz3S+QS3pf1hBLdVeBaE
SIhw0s0I1/lTO6So9yiQWuHsLcFoF8gpysAyQSGW2brsqFpjLdkUy/GCtSaDQnD/
wNPaK/vCvMxmmksueTUk4u9PwqERPxvCZs1xoZ+u72gF/f6hlL8G8rYK7dbkQeQn
8XKMCVCcfjTTpXmBJ2JIXFVOMZ0f86TWJO4Dm98m6nREkBSCtN2n7riUVHV36H4r
afc1OavolFU1wO/+pyYTYJxkpoyYrpwlmrfcxlQiuuhRtjrszflE9Z5p7oemRwkS
jO36Suene4u3rkQkXTUM56h138i2Y2ZEwrlGT7G/ZdABfzJRDTUyEN1D/uGUe0Wl
3+nC7LA10jlQMEa+0+nlFriTZPlwf9mO1LhiCPZMeHmUIU31ZQZ2MgMW3ffoDqKP
KvGSeBk91spfmf/QXUAqDHy+keoIkfktZ4BsGIhEUgRGypBBCPIgZ6WDOBwN21do
TF8pvzZUaExmJsccLMnzRyKL8mFKVWUvjnAghrsu2WOOlEphox4VvHOS6tMlajUo
Gsu60rXZD+Bp679jwY0vkuR5xP/ySdaVXHOj+NmqagxqjM3R0mrtF3pSLvU8YEtt
8qXGaSlC/Bil3BXnE47V1DW4Ui9elpjgaLmzA6/ZvqAzJ/o0zSCvHc+VAA/4hjJ5
+Ei0Q8Dw7hlj8em1qdZr2zkuv3JzqGxIjpbZy0LByMdfX3tRMwwBO2wt6mIrvc+i
BAHI8UwP+K7LsVhqYLZj9x3lkNGjY2Hk31DT67uLUVDPDOHou/OAoLIVygBfVJ8l
uK6Z03gsboBY2Uj8peJjeVHhyvMH+FXwis1dvif6Djv81R5dfpZoycRCBjUEgyIR
a8cjUR/u2ZB89lpwTTCj+N8HuJr1utXDuXyjRxqkbVT7qX2kNFkXy7e+X6zrwBL1
+N5EOOAzhoexJkeAmkWxH6Jbt9f/hd7jyik6KCveNvnPAj5MeVVzzfFMlyDdxWku
oFOw8njZlMEYub5E3lliN6y4JokeHPliXGyuwmr1BJlG0776u/ekurFGnbvKQgSR
5pRAdGUEzLwv5mwxC5SO4EiIxzkS7X2GBQdKyQP9eMX42Ztryp/lLpyOfv+UcTqI
no6Sm34FgqcoLJ8d+eC/uv5KdC/bzUuFPt9h0xKHbE5ymXWzixoA7cwbhdqMpvJf
p/auJG8dcLua18ZvSvbta7QabKHlsnCz1ziHGN9PwW+DJz/ZCEaeU7MChInkw5Te
TnCn4UOap43D99GASyOBtC3LHQ+x24oD9ePMod4cu2JfGO9WsUplJO/1Lgho+QHY
HQWRNJqr5KkPMHo9fyTVndbFl6dBZgyaJnmiCVRtVoqGHK7hDUObv0aoeFosXIQP
B6wSbvXTpB4k/15q3bJo6H1oHCWQIP05jY7RUA7CwzzvZ6t1DBEU/UbrzfDJC8lK
Cds2curvb0TIDS/+o0jUwn7Q6TFbi7a5OThVWoQf2aGyaloHPjxVAlXM6wdyJSkB
WTqQmPlcjSL49pW1r8PghwJnxrmQbZmT6GlqdpXn19Y0smpMBsKNHdU7o8A6y/oR
+KMv0eRJnLaxmO6shj8oCe1WDJ6imE7BYqbaEqgA5aHGz9sA1AglcCQy+aw4UMCt
V/VKfl0xvmj0IXj0NLhEdDX2vbhxvOWvP6/ZdRm1U9KSvHhOIbmiDSYK5Yyio+te
CqB5a9r7O5nOU8laMNKQ4SPDEOSccSXH70inQAxZmXwSHR9uGA1GUbv7zETDqpq3
vBmh+oQr6Aj3XiEFU76LddNLF2MCKRflLsf4gEY9vqG9xu3d/I3k64wSnByB0r3D
dUkq/pWqlRus/8WNzgxFWzfpol2fWlNkPw6djWogU+8ctLKyYdqD/A4APyU6OSmL
ppFw4FpbaM7erw674GPPslq7x3wzyu0wzMlgaZg20A6x2la7BkX7xkFmlTJNYfbX
zZxGgTR52ntd3CMCwbqCmMopCTNEljah0Wk+6fZWDelbm2Wuw3EgPolj3H0G6pPH
0j1TNEpVBY6aZdT/pTn99/ifkpfkfEgo0TR7tSO/id5Y0l2mwGUCcqesFaYMseVx
GGPH2sekkbt8+sMf0Vq2uiUtfpW7AawpxEEQZexP5FHd2KE61X+eZ1upLhcZxzTq
tA2jMtVmztMkFkG/dqlK//TMZBAU1hvigJ28w9/dVC8enT+3ljHkUrWP5NNiORFy
Osf8utZUX+YttVy1HLwhn9CcewkB6omU3OZTQkogGg50WHtUxBPzO2iejb/7HjSd
i/X6f4w61IqWMNvjXPwOlY43h1srwJp7593C/m3bpsfXYFPvVXw2O70mSRDBSCkK
owkA8o0AygAW/5iRXWcToFRoiq0uA1o2XoSU7ULWxmbFaYV3AEGKM8rquUTXnSIy
jbK/o8JOVJRmrZulRRpN8z9Q7T77y6ZEpn2MNNrR1+tY3HJVLz+qs1Z066klUSQH
ucVKrQtkBFu4BDvymdxMx0J6/K9TRya9ugEjUZ5YC1mExzCaPxRpETnC4khmQkOB
GTLSo0b/5yq+VlyL2ZHJ2+v1W4g7+z2+oJO1FsSCgnZozDjqfIwf4Yb/NZCbOLf+
9KN/c2QLdR5r6ZOuvvb3t/xbGo1bZYcRsLagB64pS++/2OnB7YA3o1Y/KV1ekk6L
GPngTeeUIfTEk0pjvheRkPy1dtiYHUuoNC8VgMeWEqZ3sooWOAIJXf0JX5FqzSft
QFrykOZHGAGWIQmAxigPv4bGKeyzWQ5da/GDToySsb26vK/cm1BfKjXtPjxW0KZ9
614j4CRjZ1J0xNf1X8VkCa6EB9J7r61eq/spJgdwOij+bZfYxIQtyET1cqXoB3Lf
3l/Wn0pfwsPGfzTGa4w3OpNO0p6SXngjuluKFVZ0MMbJznUv0K0Mt56Qb0fz5UMd
3pvLos8GPJu3wNeQC0kUlTUV02iENdoQDf/vAuE1H3QIeLyi5WKjLjwOKKp6L6vN
nG37lQjCC85/reUS4feDQ9DJueSCLFskYI/0ZR3Q4mAkEXe/YVfRUmvKw0OPorMT
RRUPTtuYcmpNuReYCo/4N6O1K51V4eaydd+SFPysAF79W+KTsIkCA/thr6+6JRHl
pn06c1KiopsEug7e1z1Qf596bDhOrJDnLPoV8X8yXlFXJ4xHsP+3rlDMzIEgridV
JQKRFHTEx8wpkxMd1zckiwjrxpNWvOl+RoBTtu4yvPelabNQnTa79p6/ZjWwlUg4
TCSp8UZQZSKnLOQjNdWDOTv/5vDy/j67ks69T0ytiPosSNnLPFIWpfgM9ajRu2AI
/0eRaFz48GZAcV1q+Vccnvh10fTPAlibH2D+11HcXxNy3a7HWlmTAJ+3R4Q8nPRb
FAWVkeUCUGqYUH9bi1ddncKfvIYhf/sOlDzNAZ9ySRcREUi1fCRSeh8iFQULZU5/
pt5MD8czPSK2nEj7NbJH48Tj2EMPU4JnNmigAFebkGpKdQKBLNcVvbh8/V6jWQFl
yOySzCLfp2sg17Rvphs3215wE7s3xc2aBgUAFlLZLIAI6lABNjClvvhqlNrGGU1U
5ThvldxDZ02+u1VsMZOFUGUlQef8cfaz7rESzPyvMRFCO5SZDwhBAg03WloUbTkJ
jhmKuUpWeRzo3TjCe8xlUD9sS8qW0nxOi7KbBG/dM9OL3n1IGODTCOt+G3vKNhkQ
HIA7qLm35/wyzWGHgHeC7dbR6KO+kHWMinwl/6yNSxUilcMe2mqkQV2ZIktcMytS
xiJeq+WVAd8QGkl09GwRhddYDuM54WXq0aOnvOpN75n0VVMbYf+ZKrhbEq5ZWniq
Ec9vjKWqw+IA5de+rKOp7OzYeNdL/NqgnFsX94ZTOAOKfTeTQN2SQreX6ZfU9T7r
yE/IOhCspvE1t4NjEdwLazHi4jqHqdScWNpNjKpgY/SuN8VwplmhsDRJZw0Q8kuX
N2HF41VxDLITR7oloXr78MzgTsdgxLhraSpEBONfUuxqutiLVSzhg/4GRXvpjMic
A6BSVOzVYZqN3eUx3NGoOEJpKllWhLX+VVgKOF6ssn4mUZCsO4k6EY5bJPjYZ1yH
qAz9TXcyC9yEPDHRBY6cQy2iQkeGKhrNbjaeRlJ3A02znRDhKkhgSnp9lQxBaT5/
dbnd34HK+N/zOsvmZx6wtr4DALS83G4hTdwzsHARUU1Z89ypxpeN0WfW5bPyOzXD
AfWH0wYFqsZe/KEZugSsMfgV28XcCKHees1udQHgcnIL4b5EX11FQJfwYmMY5HE/
6sRy9+NTCdETUHM4Asj8vJ5wsEoLRIr4BVWLgbVbpSF2AozUJsQFUCpdXXcedxdn
B0LJYMDxK+Y+xpRfhR+CMgDeoMyXo+NvfnO0+MRr0Xyj/Qe+7ZJAz0U51r+AGM5l
4j+LNT2qBUZFQPUt1d8uFoWgoBg+3lP+gSrj3cRIBiJId1nV7FQwZGD1Mwt68l1P
EcSgsN/V9wO/YJBkI4t/vwVy6vdt28koge/OMaXngantqRNuwhQJ5a31B9AvUiiC
KdDvoqcRyY2mKgvGxAt3hdq4f9fDv4Hi4QNF8PclA9/Vwgdgpioyr13O8WlWKw+n
DIFqxI9MUlsWmEAbbbV8Ew65ZIiaPnjVQ3QgXCp7aXl9s6cYdM4sTneYucuwvtNf
GTAK5VKYIwVqWrAvFO1tk9+Ct14tnZlofyr9WvL+Z0/Bnd50eEWx+XMMWepyto3a
JVNQXYMQ5owCmHo8ALNDhYiFUiKXQA2yMxQdj0xjINMmpyQwGHAxEptyV9b4cQOo
BmuUOM7V6hY/SoMrSduiEkmRSo7MegcSC23jM4io9Td47FUccH464jrr5KNSyS2G
iRwu5hOouzBRoEMv+Xztq3VV90i0FTXihscGHKq6xzmw2UWI4r9hJmrLXOk2y8rU
s2RhrJz6JgfM3sS4TYVp2erCiyCl+ol7TuApdbxBDXcVGrMTCyapbewqx2LkasBV
/BxLqsOKPUdx5OnZIINHM3fWSAGm1pruYsDc9VYM8CBiXsyP1NUghpy3p/7WwaQO
wbY3iZBmTyOe6oz0Gnsur/+1q66GksAyk4ClGcV9ngJGpZk8ZGjOaUMMt/Tuns/n
/VM2CK/OKGQNwJfb433qpQit9l0KmzejbLAluLUXsugToZ2QQ+uzQB4yjKpnPomo
yqJUATWhT3gzDvSrFOuAM+9E0gqxBOace1UaccC7nPJFTE0T66w8EDBL1sjAPiJ9
GAFvR9gXIt95PheRgF58Sg+5hFO4N/qyGi2Y7fKrUuWel+7+cbWkOqVW37DoiB38
+dpU7y6b9vZ4lnPrqg/Q2tiByEGdD5l1m6HoJzjkwsIEC3bCVHOs4Z5rVpTmI1T9
BrpKmmQEiD48q5aKGUVeuW9GEm8gHheTlZI2DaTSJjZ0JDGjRvsEIpTNPNQWvjI+
+Qu5tC+LB4Zi8LClbCiYSm8maRvJmtjReT1dBWNNrMQYV60qgh1eMbD5ZWpZ9Djg
0WSAQHO8WGtSkl3MXhCsT4Na7aGsvLj8BM7iobPEFHcXFzSO7gehxpiSupowhvd/
tv/MiqE+rGvTYOhkQdJcwyfMPqphLLfymI+xZeR+8CiN+nIF2F6DKSb83Yv6+IGw
wLRR5h93HiW+KUlK/qDCd5A/hdLSD1dPth0Uuekcg0Ku/k0MDeB1DUFBmqpnrUGY
YzMZSI5W0iOPYJ/lY4DtFHoe5YodjhXD7kBYzDhDWWf6j4FpH9damjajdwY81w/G
UfvC6m9H2lpDvVXI7aNvJQgyupP/Y+5abY5a9Z02U2JvywfEZ8PJfBvXfULgk3bo
JJ29xKvP9exsxAny2gAGU3fTtgaFGrAnwhRpmWvd3XyWifghpsVfV6EZ+iJCzxoh
47CSY3qgtY0nZPKh/nKoaHqHJB5Z5JC53lcETwUzm7yHaOCiDM3LyBuPjEQ8P2JG
9cu9SXKffqHJsYu2AI/7ACconom2j9/aAsriBAIOygWTunoXU2LKCKpUdCluIiQE
9hNv7lyDl/2VGxvxw08FHmH5p+ojy1K08osWltGoXOKeuzYxaK5eav7rJMV30610
c+7tk7kPJZ3gUgSnhDOG1lfIYax9HdaosGr9Z9MwQzrue1WddJaoMudLkijrQbDO
GEKekTA5qEXCjChoVmjMUReq+CJoXJReJuPBmeQNllhuktM8QUXFfUIl2AEavHFJ
FRNzB66LO4E1BWZK9GD7v1ISFYJrnxcSfENWFUijBoaILmWF6K3jTPC575UukrzO
0p86r/AgsOKmmx472bSWbLUdHtitIAhypQrARWVsTg+bMDBTFPm8XAYhmKYKkrQ/
8Z907yRgiV4njCZ/V9bDabS825pgmFsLthTIqhdN7lhg1HHh8gm9fJnRYgv2boGc
CC5JRtfx01+ebGXDOQoBXZK+IJjmy+HBZgwOWjJl7Y7sn0J461fRzYGatZq9DHY2
VarEcq4L82GBB0e5/oY3FUPTwjmXU4fHTryfzbilCCAlqfCxLAUCsEt0TZk2jcjx
SdoN3Zr5FzGZgx1je9jP8eZ4VwZsbYRB0DwWpMGmUwhNdxOByL2/aSERMQkH3fpC
Od9LbR8Pvfp3LNUcBKSDZCn6i30InF+cZrrGOw4oxsZfgw2gYAWHim/W6ckYOquu
cZtG1z85qbWyNRcnnD2ZRAIqCS3pdLnsALEJwtrWC115uyhadHauwP03bNd/D3c/
5Et1GUV66TEYViC7KGiILP6L/Cj5Gt6lcfQzxuQUBUBg5Ie3B7oIWN9VGxNHyuqs
VcFqeBh8hoiJ6XT+xeToAWeX/AThIT/BO/0Z2FhgA/U391jHxPeYzy1yL9LPWPM1
QZgvxhWeAN56tDfrCd+qYAEGp+WUt709qqXGVz58DEj9q7eW5opICSloNpYXGn+4
DetD8lWASvgY9JoemufVkm7+bHS1+XtiM8yExmeK/O3+UTUtDB308Zw+zD5i37NT
ir+GvHJY5+xIbefS4I8+yNkyogqbzxwfh04Firpx2JmoINyYnq4v8Jhr0YHP27ZA
XSJ+nep3Wsv8veIIy/x46irItO40Qo71SVooX6i2ZDuCCn8RUgkC3JyhILjFraxt
XqWmWdKKEhVRHpr1L9Y/1tKKBcoFeX6zamLsANIBrkGW0GKOq/wTu6Msf3sNPK5v
BM6BBWR+ZNcensXQKx3RldOK8jDnuO8arNQRb5RWrS13PsdZqkAJW1VtYH5s/sZ3
z7OFlAQi5E9wrcaVUmIsR5/wpX6nwKR9Y4vywyfBe3fG1okWfM2pi4pIynH7PW6L
FITtK54/DhrrIPZxSpMaIXkdJ3aHwgQF2VlouM7TSMUHxMELUOH0icJzdSN/zC8y
3Z42LChh8Ys+WUqLBndt3Rmn349qfA8NWZwpsCYIj7BDTDDBuqVHQMvSC+x6Qt03
goCdWNwcpmrP+HYuWy/uzajYIeIe4mEQWwVupLJujj/+wh4WKHYib/upRoFyArxE
/YPhKnK0J4nFxkPkrJZSAt7ttrUPw+FdA5WromVzX5SAYG9lRMeNwoXH7bIb08bC
zLoXsAFYBzbTgjjv+EIPnEvqoDB69Iz9IzAZDbmmYvOSGF/yoQT/Bhr9RxxTx2bi
asmwQV41Z4sbjubCnUl4qksvxzg+2dVZU//wTkAx6YhYJvyNXsRLqzmI6FEIpG/y
w8sH36LqYKKfvSXPrisxSIQnShs/MyrULkzZnCPO6UA2ifgsj5LqI6U8rvxx2xpo
Tny8nzL7mhd+qCSMyd0Kx8uVs0Uf5g36M5Riwu78komDR1jI4mzP2SNPwVtaVN3N
r/O9bivoief2AU2h2LPwy4LdphI3WQd27P1bcj8AI/+UKTTsBGQ+ISAIusg2vTZ6
VPar/ydDIJr7EXGIOv5EbOMSVZI/DtIN8RFobdEedMP/PaMe6U5RNdyGkz87XM8Z
QkDeS+d9kA/OxDPBj/8FJPWo71iIBKNCRCHRrD9sKSSQdVGbkJV0krPvGUCZmW0+
E0CQ0fOGaSo5jVVXEZHxz1+0V9e33I3X1DJHjy8WL754I+mJe0mENYEn1g8PZGVP
oOPvdv4k11GhqXqr5epIKAwqno4iTP3bXXumgVCM3B3IseQpDRiD1mzMHoqx1Fdk
E081Ut3klxPR1mkHQFEpx/XveaGd+MN3FrelGwlR8CJr6wHvs6cOT/8Z56QlQiTa
v+H5IN2F/xapeuCWbGTmogq7fzXhvNobvqXgrSB6yo/lUTOLLpVIzT8+FPiOGoaH
XiXIu8JQxGFVKkzGZR4FdLSc+Ju2AvFNd2jUnxyjZ5mv+7Htm+GKlqSzPacKJXad
/QhD/j94b5vJ1E/RX8h14Cmbx9JFWqj9Kw+qdvsLvGBwXyA98yR1tkidDBNpgf1C
udDpgwLDwoovU4rHrA+bipeNe5BRwYWM7ixcJuoAf0+S3dWRQo24Nbt+fjvO7OmR
NdBxj/1Fn48MiBajZxPJSy1Kh0DQCn5hIjyvWx7fyj6zUn2AKQ74idPKYawxFbUF
qWVD6TrjfL5y1jNYpyTtRZumK+W4OclX2DckvoL7m7gMcZvrjHVmFU1liPE4N2t+
f1IPn+n5Czw9ZOefaxI2p9YR3knh9Cajfri1BFB2JddZSgh69Aw0pQdJCzp0F5bE
EOGS42NaIo5RmNrgVsDR3l7SdsJjMoVrJmhStpZXAkvcGXexfaQ/DDR0b8GqPAAg
VOwQkra1XRER8G50zOo9pBwfXbYF4/XbV3Zlsus9c+viuXZ0U4d2FkPI6VJ64rCp
wuDeHIdOOmqPoXSvesZQi90OYqhuQJkHDSvfywSTbVaGi66UVLzSNFad+u3lafHT
JwwYjRHelPY6k2k4AUjW5Q+L379Ua/0VgYwYkrcRwUx3Co+eOd2Bgb3m8DowEF8Z
BNkLJ7Y1ixsY72zZLWycHKT42EKpoOOamgMTkawVgWMnaIu4k9vup8h+xu4GP5mr
7VA4wWKpKD7koHuaN9BNfWUGM45HccDpoa1B42b+Dk321Z/OsnWun9Ak9UWm2DfT
ZaJzq69xHncSBhpMgEhWw0jqMScMneSiX8dtTQIAUHW7EGqCw4/8Z57lnfP3tpLm
epFn+ocZftTYThUhD0NprCUp9dSUc5M9QRcpgq5P0o1LyVdAFABaAFsxK/bU3HlK
RELsZ2AXaZopk42ZQaPC4xsAPhLn4SyJ1vTzOodle5/gSpnBhnUY7GXky5nOeOqV
nJWSSbv4+GbBAwHiECKKojLCPlKVGLtqwSeWvmVdRb7/+Upl9LqmpNnS2EwxzJ0D
MSk+qFrNQ8ufEcRzPawU70iiS5n5a6qUObHSOen9bvemAbaaWiyBRv+GwcbL9AIC
81njRLzBfUOaZgtemuU8sOmfS5DuR0XsBJjPM3wChvnTEexzHdIgvFNEzKr+3vAT
+81VVAfbzIaY1fPNT+nHraXbbmGPwpIVnfL00H+JRIZh5V1A8I+BA4FLB4OubpB6
2trtSgJeY65T01CK43XcWXVNAqTF1232FUcM8dyJNwBQQpOl4NqgWqZkOdJDHWLd
FkJRji7S29ishC9RYMhnO0K88GDftIPLy3OnVtHyIbpRGL1MY2GcWHCCMOB0ORZn
y9YFUe9uezcecPPrOj9N7eCO/JQgCsS+hjp5ymTZ9EtZxzZf9mhdFRyTYmeSqUig
ziZ7V8fnkOnpnoHMwBjQTyNErOxOmR+QdRAqMu8UYAk9dngT3bS8UltbsMJLsBNt
gv5JqJcf9lRG6qYuLQFCM3OjdiywTkZuwgSFSh7bNm52LPGYI9mrREnJSrarDWYp
dk9ZFvzSp/PW3U1OhtZwhj+BnEopYO89VCXEREwB5r8rwre2LiQAcLRrSZdlsQDy
0O8bxq3W3QVWQ3Q2V8imwZDzdhzsCActmYZDX5GX7uviPENy6l8qZagMqt0dZYQw
bvetMi9G9IHoL1+40NIMYH6m2vGX1uO2jLBCNB6BUq4D8lRIwHuAdR5g75XX2qJN
o1XzbV64o2Qyz2OANtzX7P6WuKcPgMvAk+12gZXpohV0ksdQ6DnQNghhhG+/rz64
xOu4nAYym10fw46UGWzmwjLHoTF9f0qaWPy+igU6Uq+pIaFrc7TOX0y/KiU4vuWY
ChAlpeZsmPm3hM4HTgfIwNsqcTIXF1MD1RiBc0e/xpB/lakqtc9P+kvgoj6xS3Sl
Ri+UCY7ovjIRGq44VPTlyRmat94j/U6FVkF/vusYU8/WvGc69Qizef6Axy21SJDL
zZzngN1Nsq3tsK8nHSj6u3SidGgDpUPFW1KGZoXYbhj5v263MDxBiAuQMohpprDq
EVjK2ax6BZc7HEnk5mRtmpmVF74vD8vMOHKBPlajMoyGbwMOgukirPUyFdWqyP26
iUw4Oywr4byjRy350VadfqZUHhm6L8OUKdNv3VL1PRT+aE9XuacdHu6KenjLzATt
dCjT9xlTIyb87wxEwrQyuqo7lJ+BphkjFGxE8s7JFAad1pfYJXhAqOxc3OAnxDYo
htIsfQpfc151HGVEBIjxTw4KTcHBmcnmVdHPKgVqNLNUQaEM66KV0vq3L3ohey2J
HPV+nz+Txg2tLPZ9nhR1b6G/HQTdt1xT2s59ID/VdlkfU17A8E4qgfjDL/NxLru8
LV+BVfWgKeyHwxoBay8mI/zSJFq0vtRTaBkYkTzV2/8+mmdtgE7FnWB1Yj3Na7CI
os/4qQHxJP+TbdiMRNcCaKrGyFP3QomlrGSPbj4qKIo5pAzBpyX4hVwlXKabvo+P
yLFSeH/4zOilwRpElVrE7qQwIMEuORDISiT1HN7bAOPGCUANKUcGjgxN63Coy7gi
EvibPXUkx4POLKRmglkrVJs8cQ0yvS18ln37ajorFBxTidNziFakcUohHspmkqmA
cB+YrAdRK6hsqBT8iVjf9U5CJh9n/Z+IhexS6lrgqCXptm9AlR+KV84T19OAYs7X
HdEyovWTrb5n/5kayfpOnc2bAsZdiSiKmP+Odrpvu9VS2fZHitdFRykfzHfoCv7U
i03sp9+W3JmpAunpmEqxqP45TUTG8RK7OG7ebkhjsPkiAc343HquMvzI6OrDutWS
UWWn6xJ8KrtVR6plJnfOEIeZ1qVy4US5IPsazrKMdEz6Zls2Q2S3kNnIJ7voFAtx
GTm7WzbC2f4vfqCmOrWPkjcusvulZEwKovQPWVGlH9NiJaO1NHSWgU9iYJZ8T0Ig
Iwr1b9O1LADjc+a4nS+v4DPT/wrAR3ArMeZZWOWy28p7K12TX/cZdEwMeHklXnLR
yFDdspv9CgsUd55dDJ4HP8gXA+vqbUie6pQfF5nOmfd+AtaU70vpIV0aBTf99tiW
kyvLWbglDvLezsAeqxhac25CbWzivEFjFNEAIPJoXaU5oielgdUwFFpdABJ5Gh9J
jerfCpek7nKHnWQMzEYb+08pK3dn0bjUdjBb2N/KgKw/q1NvT/GJBEPaR15OnUnW
/vKAjbNXwx8QAvC1V3kMcT6xdHde9z90YR04f7R2EYR/Wi2o1EpDVj4UIgAtpL55
OOuhROVc3p7We1e5w4s3mNzrUgwemOGqRkRsK2rURhQxrIalYTWe+HbvXcR4uJom
r+hQwPcCswRuwrkOfgy935SkIwn+dBeKDG0fxuj3GLuuRi+MwVPWLtSszvcaJ+tf
3pERY2py+YlUI8D5FAzSdraBFhIappjNe6tzvFrmkePI9K4A5ycbEct4Tpq0JMBC
qQxvb0KCZPdMUnktMp4y4XNyA3RGevwLIOGMUV1ii7h5b+iqg1WC2UAoOZ2s+l/C
S1C0fzG2dQmQ/SiRTcueQqLpgIpJANYOoQNcHJjNP+QUp/WCMxNH+wJ6jwYyOIDN
7mdtnP/kIrMuRuR3aZpSuhtGIYunRk5giv1/jFNeBl/SwxfwMl2HY8EZ1or693EP
w0ISo9BtitKqn2iReYiiMVUTO7tm1e+NLK2m9qlyMIHVFbmApopZgsWRNL+fNxsF
FUiN05NLzQ8yC6DdEEkaXtZ7tq/DpnW+3aI+U6YX3T3iFb3tX60Rt0CI+yB/DMdL
Kp6gNzyn+9InPwbUjW4OlX6MlP022PYINiwfUUdqY/zlEFxlNx1VfJspFcy2P7g8
QN6o8lpwwRXG9i/Re3uQYJz7wTrRfTsLmQWy+Ev4+f+i6kSTDxaWhTpGjY2n8Wni
X0+XcSIdRAzT2VRjOUCsHthCK+8S3flGHWen2eKsxePpF0dNfwHvZyhGInBL3MyB
okL2cqnp72jkr5wRM0W9rJshw4SY8FhHFoNgfnQp8gaeke6Q2ED4KZPOvtfIv7Gf
4Ef1xXDkKCJQJFqshPWJQm9XL5+9TCo0Gt8hNXIqtNJRg9uUG9EEhh6e/wZvjsU9
TtATxM19n588vugVF4nHhL9yb7FKdaPg7bYIaLg4TdfwzBzQMtUWzoT22fzjM8zh
g1/3yvbPMjdm8ROU6AfxvTFUNVBNbyyIZMfmimVtSvbu8jBHNE6b9Usg0ZxUruNN
zg6E6y6ErUY9GEhCcPKvFWiIqN7Cm8dJCPrjPeJVrUYZxXaB+vw+V93Q58qM/g11
/hGywu4T6ShB6Vd/8qsp1xoSAEZmJilO+9f4QA6S/mVft+z6jjfl2CUcJNvxrY42
MOqTxHRUMDUSSAneW0Wln4Y/3rkgWckhcgZ3fI0+qfGeIkx8XKQMkYDav/YbJcJF
z3GKNtCdrTXkil6LPgS9miMaBClPeXx3L4ckUV6Bn/2eybJLaU9+hoZBz79DC+Em
5BzOf5jN+9v2BaJO9J6lGazByQ5upSiIm8SmAVdgznoHndQaGqxPLNyt2WT3UtUU
9Jo1JjaNOVuT8GB3eg+i9xItxFBlzWDzS38ABXON3RMqJqjq7P+/H42bbQQ1fb9Q
Exk/DziZ+G3yHA3RobkU6bsQb9CbIs34Cw5o8tH62TCvVtKg/J30RwQh/h7Lebpt
RcfrWpWpWHOAgE0UF23fr4a4co2F1ghm9qxJjmN2jdqi+Q2/Rac3MiWco56PrTZo
oqO6JGgtYuYVwnPOBxVLGPw7NOmRINIff+YFY28UfMcgOS+P6G+gJSPHtqxh7C4i
aEzEo0/n98gdCulqQtn1r6pwTPRvTxjdIh8rPPUVHx+wTq4+btWQAUjrJw717H3L
AGCTI80Tm8I37z62BUmnmeI6Z92XLP9Yy4qzwqVJVrYTIN+PpwDlThs9FHvObz6G
E7V8ILl/ldZ5v0ExYappgV49HOPdwdE9Rk/iPhJ0v/lUeL4t4LVqXMG9WKLumxq6
f0dw87uIw+l4HuvtCdYpANmeN9c2YCS3JjDeXsQdqvAdVXB8/Uxq/R48jLnHNh3w
Xkjf1bNH2F+dMXQOWgbLGMAKUftHyZ5B6j3bA8gIlhs2scVj4bpW0oLpl5iVLJtS
bDvF8PMPl9pIceMrsR0DoJwSP/Mrx+3xsiWY8tH+i1Wa74K/apfZVpsHIkuh1mhq
DT5bHuIJSlJpGEwoHX+86vdnbLelAC4JXqt6nn1Tdpqp2iQv+XF5Z4L6+Z9uxbYh
ziSJ5QszmKXn7IV4aNv82W0b6bam1oJ5LBope8xOFcmXe6YW/f42nl2qHxIQjpJn
8LxYFNsEdDQzKNV5TxUFbqjKji0uHInuGol8tBoVXmelO6XGh16BzY3jFtxPR/HX
QSCV8QsOKVa9sN/MzHg2q1zcPiTuW7yO9PJbowjfXzzGGS3aqiW6vpH97c1x7ZBs
wPkcpYmu0qkUM0TXFmZ/jJzczf3gKkGS/5e9ljvUr27PQoSbi8EJAaJgE6MaE0wc
MqOEagse1Fj0y/mFHwGC42chWVFFUByTBPpZKcDokPo4W3pcY2JGPCVUBxxA6HyZ
nHM6870TV4nyDW1tRAL4VGLuBIlj+Pdv1c2ORW9L4YsdNi5MPRXgM3xdkjduX8EM
NQ+m5gcck6pyuzMB5T8EipKQwuNPXB6PRA0wS31Wn2U3Ayvf7IgfmXzq/oABs4uv
o3CUz+c6RfRUdC8D16I/xW05RN7MUhtSXE7MLOnEo143ruc5fk1jPm29lBHVaZuh
C8iTuJyHVgdNCEizAk2NGiUo3qBtYQmFspP+VLfdL2k1t0d6aJ+clFSQfeLzySEp
oLgpKP+M4zTT4XOuc0GCKHESGiE6AxaywfnWmCRJcu94R48Jeeg62Dc24UEY/eB+
5Yi701vl6BXoUxPG1kfFp3MZWuOCl/FKvVSC8QxJtmljtzVMi1uYa5j9BO0STO9c
XcMALfThC+VLMnT1Y+2llEibL3zTHA8rn3DyblxU02kwJZl/TJGxZtTgMIqzoIx2
TzlKr0H13BCDmdfFGpHI2lik++aXgdnSnN4sq6JeZwz7sAkh95ILROLlmKk9KeSQ
LjcLNEda6damX/P5ehwHtawJ80t8JwWcz1zT3VLQUZDQrl4mjLyMZPRT/NzQf7Oy
N898yg4OZV8mtDelBjvRf/l+jtE9SuyTbj/KY87ppefNxeVfUU+VodPmrql3YHvf
S5WhrLVKDIvwHrMfFIhj/QqXd6MLt0sNnnjvVXn0CehPsnHUcZZzvcoh9CsoyGdc
xRm3y/z77zzVuVp/qJR6eiXUz8/SGOVG6nhKqK7Gdx43m/4MNHePSmtImoM6A1U7
UghmsAOii3sraNlMaWE2lMc30wMypIqfq6FFeumWMIASssJmryamcrt0ZNRW+d0M
R8AHU5dKdqgkBsjDwzvK8qcEvK/0iq8DxrokCf65BJijXPpaefwLxp44WCm65Qcw
GQXuGmIm9p9Akj1y6PiXwBGiMt/GbsfczgBDRmCTV8embalzKWXXTx3AarvOEu1e
+IGa8GWaROtOdKiYw9vrciWWJ7mIyBeb105o65RZeA1IRXIFqw6mhWHCcVI6Ne3k
s8/bNBBjdtWhWndN4LdY6dCYS2f5LNUjowtFpTojzBMcC+rkii5EtJcdYC8bI8nV
unOnJ+lxjsizCEHiuzeu4Vo0Pln2TzyeRRT8NdFfJffrsG86FSXO2Mn+2guLqLkN
6K1AaasW6wEDre0FAr3DhZbvBefPLkxkIDWk56+gbLYpHSJuiOuIWbtkuVIcmEul
lKyX2lAF6G9e98sHPPFhHlmEDwy1CbvwLjQympKe5EcEzS3RqXexg+NE86GvHJfv
XMtDxA4EC0KpYeogq7FSEwVIQ68bRk7vGnDOrWN658LO5Vhra/b9DMPHeBBZAl8J
SbeT/UcjPmWeFZ7v3aGs+FYjUyBeniINNNIyQDSfjJilswKyVLAYoRyKW2hwrlMx
zjFItGG510GA0iyl7dP4X4+LN3JxLxML9OijK8Go1sR5VqksJ/c2bLfW6McdtY6w
SJA0SN3SaM94Y3YnPwFwU+Nnm055thq+2ean5s/sgWNVRTZhNftTSNaPqsLE7rui
MnQgu7smCXgwSWn1vqAAl/Xxk83bbEF/IFor1Kvc7wkn1KvcGt2qWj4XEGT1IsVq
1lmir9wRch5GzXk3QOoua7xbeSKZcHaWMoy1rM51BYyIH6ldlW7D5nO3LdSOX1zK
1Ff9CIgm6UVuba8PTOVVryAmYI6ewNV8oL/NN29HLLhd9lEIjoN9jqpgbOpKiQns
cs8vZU56H+XavDmRXjYU0OHOH3OLzOKb8QwocuxyTxjeI5Qj4+0IKSkNwpYELwwh
EPt6OzI8lEw6HtX6QheZc2pYXj/mCmNu4+/4XrwNvnc4b63KGouCIOjdbji5SfVY
OJ8PWLRsupM12EBx1XVVvh4FoqGfhOG/Ztdy8sG/DMem2fJj9wJVEvSupt1MPYoE
OZx6+67xZt6MqdLnEkeKIGgLsIENdqM9i1RKks9CCBj3P4rPLAlmJzjBHFRXM/aO
Cl0HPMP4ExkxfESuhxUjjwwzNyijW2VhuWXQp2juCbR+LLkHK4Nyhwt8z6ZlIaua
38kFO4cVDfSCM0QczP+V5+z3EEpSp22aM7Rd81k43y/GpLBaWJI0EeMEMf3R4y1+
1gv+q3sZdz2mu1wQPQjbrEJVmZlnArQsKKB7b8QqXpqPAG3iS2TPmRVtJjcnqHRn
kSBISsV4XWMczDBvoW91jIR6tvXMTUrwzAcuRpK0ea6njPrM0hAmdeWaM1BAP12F
1Nc2yEPqmgbCAIBOBsSUcU9sd8vqXRKZ+beRfz5qArLOQsFBYBrLkB1DXn248rCV
gfmvRnLi+0lDybqylTY2ahO1TgYGN87rqiSkSMCnZeiTcFIOtsHPnphooJP2EfKI
rihFHqcdTHhbvkEKeETyW8xlUm+njHlzjY48u2xOZO/tsxfy9hfjIivNB/vMt+TS
WlgdU2UJpNpbCwGN0Qpm/6WBztiibKlI2yneSrdQJbodRrty86gKuZLG1M5Q6vs4
oIgt2rxc+SNVXWgGoJeOrm7p9APbp7ZNYHgj1y607EIo24I9vwD7g+64w9rbXwm8
fC0S6m+TNUUgEzFelIUifQeFHpiU5mOkDeah4vMcR/MwPZEtugx9BpVcBqglV7nG
rk5+bVm4/XM2aVWRiYdk23ab5pvHxptqWf5/QDE6EUWzjeB8lGEcqY/e5VeUW6up
4tBOkJlruVW37jxgqfFvD0OXkNv9gPWBneIYmAZXhRjywvqijw3YIXqPG+6a22Oo
T/pk6WeywKiFB+QT9zLUArwTrL0jCqGOMbAWP8JgotipVsMlFls77g3uODOqrtsx
DAvZcrZdxgpXgNpCyW6AlLXvxdd/djGY7KalKZLayMET2ETuthbJODd3h6B/kgyj
r82UYw4P7QEfrJYJAymTKcxsItbS46fI1NIkW+PqoZEWfrk9iJU+zyP7enJDMSTg
qZIRwOfyuUZBD//rPrsxbJMjtF5WwF6RNSuu5FPeGi0m3VIFRvAE1LdrdMGBrDig
nXwYMKej2yO4dlDJ/Ax1ylVVc49wTAUEuYchDLipPl+sxynVWpaFFr4f611OiYwb
XJJzXsSiuyi3UQLJdCVsM+6I2LkmsczzWYJ2TQghGquldh3fp4Gy748COVY/3mZQ
LGfnQMqAMUxqksXUk7HcRUVhVNx6ilkH2XyReu0dpcsJBQWgC0tZZtFe2nCu1czx
yGQaLHPpcZw+LIWFVhAI8vOztIoXfkymNhw2krIrO+omzrAv6m/z3MGmPTCvdRBA
nb+693Cz5TBGzIoQPlQhk3G0X05qlprC0Q2XMZlWvko8LmvDuP508xq72LWL35zk
Upv0ovENrw1QLx/impObMpTT5ohyn45hQ5l83rM63tLQW9ft8/WZTO9kdxWoW9vR
LCyY4kCCvmRtJ3U6pmjPzJnl1WWbwPItv4lPjSQ3W+d5jvP7Cavg1j5kq5x7YNgi
9tdXS9PuA7VPi2yweW6qTGPDHh12yHmbVurBKSelYGTKmF6mpOJoJevALaC5zj1j
CpwQFDE4RGCNDpTdKUt5DGWIoYZirlUsZw6VnSxOmy6Yl2qEJJ2gwGVjLwUpexT5
dF5pfm+UEh+rGHOdsW04z5Omz8J9UFrOWwQk3OOJkZP9kt7ch+KZ3wmXQRAkbkng
fl3ak8oYA43Ln5JwA9Ht71HoPLyQbGSElw8yStuRQfmQyrT0ZCTn1+/3AymIUA9v
HiNu1pW9hQ55VIFR0jUA9PR3oglGUvynmX8qvxoc4h2QGp/hiEcnKkBUM3BCE3nK
Drw9vKCLN2/qSTv+ZrbDFfPPfpOnV7e52x8uTHZ5k9Dwxx/7K/bHgFKPNg/ne8KI
FPa2+lWuOCVVCSsBaDdytFvtCrjWR9JWi2PHcu4UhY8ZIGiVPO7ZdpiOHyFfiTdf
YHk6cGoIJwNCcQUSz28YNv6BtgB2KJ94gfRdJdgHXO2nC3nnuZX5hpJy1yKfDWKx
tW5CtT2fZXePJqnsc/FW2jhSTMlHcw/DAZrD68z0BQuyxljJoPDNwqQmTQ6tZY/B
cfASNaI+sntX5sHJ1HPmboV4vsF37+/abJmaj2rjIgjB7WnmH/J2ADZNjegEsFsj
a/7BDtHO9pcLTn6/hbyzh0tVTNap3LAGxYxLf4Lb40Y4/fg5OJ3bEkOfdg9iCS7P
WV1FsB+nKliRK1To0QfXCoweVwt09XWDZzPl8xZclG+FrFsSwACQiilw1hXBuH5z
AzWFWkpmwCsO0Seq5iU33vdH6cjFkzEiJ4XPgLFL2MoxKFDiiptUptuRZhgW6ZHa
FLSRVh+WTrbJjwFFItkULF9EE171R4YHw1z/oKpWWaqNFgP+LXpYWv4IUMKy2Rpo
zFnCPpfeYmJhVNuWTXxLq9itkM5MfNtIheqYYrLlY1pWYGQmBL2ZBFsG16/obsnp
I2VtKe5u8cR3/d2COC9HiQwVECesKb4nA39in3TaHec8UNX9cQs0/R9+vgHl7KtL
gWOOgar0cjBZRsn6cmdyQjHyOTWYtsEMF33Uk2GRw/Z6q0OPvzZdFjGm4nHRP/zJ
GjnVtL9sgvxCS9JgQuRLcl9/dbc/fJWu1INGgpJEnXwWSwgvDe/MF/+hkxa8MNeA
zyKi+n696ITTCWvzMxDpETWzjLxwVM+rxhDQ878HpQExqnDX7pIyXl4I8TaWt3Ho
VMxQl5AZK3A1Kzn22mnAgCl0Q5pN6tvmj/a/v+gpcYbLN5m8jfTNw2Ms7gRREaF7
LpytqWlkOOdDNwJxve+7Zi6eAUEV+vYt4tkoIQnEodFw/XWPXblSBGxOS+82qbWF
oI34+L31qnQw7uMesiAZWJol68aHCzTRalj5ehdc9UCiW0Fp4mCaBbHkpTdufDSB
o+2yt9UhhxHSI3ESZsy451c99XsctaI/iWXmnmmSKuFcbQ/8VxWPKbyHWzi8ap27
Zzgy+eyPrC6+hnWkhnxo/cc38/6WEBJJvISeY1HFsa5+IK/R0BaVw65HYVMkIg3/
gMlfFUNwoLT1TlOxare/cjg3nyCls+9ao/+6F73MNJsIQhkpz/7AuKfVnH4q9MqS
YRnexVsKEkQUQ6uX1L0UbUS7WerJ2NREP6HT/cN57ztiAfq+KlTUa3r17TyALo0k
6uJWoYCoz1MYvJbaXIAnT5jFrmtq9q/uHVwwAnONi/nzN6K10LQwwlPxLdhlypHb
vLGT358GikYGxsT7ZE1JiForuJZblopasKyC7oJ5bqZClxwcuwoopDLeC6mmqWiE
wt6ckWEl3iEk/EAy1Yb8tsEeb1UYqRLbldwrHwubx/+olLGAoyiVj9TugFundcP1
N6S0VkjPjVr+iPRGrvFxNWQQE9l8d5h3qjZsO7Ue3WO9BU/zLjjCm97b36a88Rmt
riguJ02iTzNL9OmxBT7gr+CZ3w0JBZtUQQWfnvi+vXWStBEoF9tz+/DC2sd6KSIN
Qcg5Dh8YUbwEluOFjIBFRBeIO7ElLqQQWg1VWt+qTnmaNGEFgTo1/gXRoMnzFLpt
BijG9Y8HvOh965dAp4OG3yqbdGULmSboT75cdVGdw5wUIGaHtK7jQLLeuyp4Nt49
bYRP97EJ7K0cdtbukrczoWkB+qX3E1KxudX7gC1g5F9cfN59J/JPsMwEzYHeEw/M
51zVmPsHIixceLzTFxEQw+hwWZ3vLIJntqYSDXomXa8U8OljOmfeX7qQHyLdPaiU
SgPcaCm6lR/d+vRzeNd/80Yx/9YiIHdbRXjFGhvsaHvmB6gor/ikhJd/UH2YTZVF
CUuSsDihsrSBGGoLBFgdP/SPzsS8R1oTSqybHaZOC323WIdQw+qE1NAIbIyAw5PB
Xgh8hT2+6zXVXb+GlB8jTs8a3588CHwTNwIJw0dHuKOnmoyYkFZFfx5QyMXNoofb
0kNIsNLq87r/JJxAEYxSkKNvtNwXysxJvfOOQzT9Pr/wVpKwNQPDy5qXrIny1u61
tqyyeOEsWJvic56ZPHLImwsN0EiEs87ViNVenRQZHlsbGpXI5v2tmalO+AuRaK0s
cQGDACvdxZDpCCLwwi1Ejei+YKkL5iWdLURI/4uK8ZqFvH5RHUuI13GvzGsoxIHH
+PoLw+f9FQB0desDI7NG/GcmQDf7+EvfvTveBLZCbeWo8jKvpzTmg9UE8dSGEv7s
bM50kUUrIzaX2r1dKW+UbIo3TU+3L6FZ8YCDET3QYjc7gbMrvMCmA0TIIMPSGxRV
JCKd8giL3tYaq/Hd4Zqx1Lc4X0RRA0hVMJrVkeoyW0L6whAk8E04e+PL5bfOcuw5
/+++MNeBbXUAfRtz7dZbgScgn9j3pNwf47Vo+QTzI01j8tCdivSuYqVghap9zivi
YAayXJswzXGqHkDCrfLTsY5umZutEPuSsD2rNnmL9X6sN2PqdagtyzCL16tSsFZQ
k6lfEGwKhfsrs/vnFnqKG1q4wMQzw7lls94R9nEgG3DlVnUVXYi0uEN/gT+Yy+8J
4IL0aAujijStVDicLzbkv9LdSObu14xxtTfbhEEZ+z4o/D9SfcRSpEqqhw2ahwBZ
3nac/+0+Im8z6oYPameD4mhfF6TTfKCnhRZH+mLWqy1GYt+u4MJkCFrYz7xPg6MW
fWp93r8tuV0HWaUJ3DeL906nbtTTvSM45RuMyuQ2zAoEA8QzrhmIK7b5aVkmZ3Jx
2d3Oo9pVmaIhA7xZu0fA4tq2MqCQlGrAfXn8RPgJXHYZoaZGIPpmOzcPGvugGkta
js1Dsaw0dLyxQsXHbe63CKhBheQdo+CkyhKzFAlfr24jLc8D1uiUNbbya8pBR0OT
nPNqmo/1SAX54a+NgUdgyzTIeiUUxT4fx89UnQuPkPbJEbyTC/YqaHivAPMhq1YU
pCt6lFogi9sFsiLUBA/bBXltj+qZKy7fe66U4FSgfUldcQfS8fFGpUS90qx4DqT1
UfMa0dlUNrJQ/ssvUzIY68Mg7Cb+K5HCsF8bneh4xs4n4dtDzCfhpAfKxlii6owX
7WFvxEPWiMTYOl/IcCPYXJqpFkq+kTLmZqak2ucmze8hs1RB/RDvm/2O/7cDlran
ZuUMDDkhPmlBzCnFicQXCudT3oeoF8kA3C6U2QAv8Nni9tiKa6jjael9cY7aiS4F
8Z1IY+p4Jpu4ZddC1Sm2T66tqM9a+nV53/XiF+RZQmWcPpDhdqjgYCT2USEhBeLO
7A8j8bqjTGt/z6X8SmZlmJV28KZZuNqCjl7LipoDQO9oxjAa5sNWF84KqL3iTp/i
3YrIAruDV7BItJjKeAVwPbM2Av6As2A+gj/VXqoYRZtgyOWYKMHpPYDKzZDGwYm+
QOCa4XCf0TTdbeLcgUmkavUzaoazQCQFo2snSoaia+Yc/YCPXtbsTU/Ij8TuFbnT
43txrokvcujlXC+NhC6DqA751yAseZKF2MfO91exb1FxwbzY3snlw63dku+bEKpT
R3lDbFpxvsM/cCdFmIIW0MD6bpkerKzglTRTUcnW9p9sYaw7SWtHBc5Mgr3/+R9m
16EzRPxQJSHgyzFcGprR366g6Lfh0zbqRjAJC+QjajP6G4KUtD5DTN7ZrXBWPbos
JSzesWFpuUaPVIwHm3L6ONwTibMdQfKEg2I/hmj3KeZsaUpm+zI3qfMqMptyq9j/
DzdQ9saqwlssKjfh3kc15ZjcuMVFIiIu/KnEsDWDEjyuMmi+hIulxrt3gdcSJv5f
xJ7nGsYyhdnAnRNTOjacFN91rxcZoENOiO3fmpBHXFvg/0Jf9FCTuoJqWMDp7KoG
IxMm/s6nI+WoOxtRG8LhQGBdpg524hpIAA2wH0a6w/lt9dKomU+HlgAVuHBaozg0
Qijh+awTQnBI4+Q7QGKVstj/T5EDD98BkfAYk75Yt/r2mMByTPdTrxRalYoCU6nr
OaCAN4YldDBI+3WpNb+qxIwavvm1T8LHRBEZYwYEElUl4LzLsgC7uhaC0L3npAAv
LYQ9ZKGhIpAaICiCaXr4KYTbAmPVOFpf2ktYtBj6/bAPUVm5F9R5H7Iuh+LsIhF3
cPe3dCCqnaD1Lix3sNFqhx0WSr2KS8Y+PObJybaBavebrsXOWfube662h/s0lH34
LicTKVFNzaQc4ZaAxlrs5V7LTXnolkCBtnrzZcldWFxB12N+tT/16djs2X5JFmeg
lbO5T89mGwMvjXmyTNI26rIZVK+BqVhjxrnDKeLl1V7hm8qXD0lm+M6TDkCLDf9/
8sOxNlNS7eCWI11AdRuD7KRXnZ1rpR1y8brPm09APFN9rEWyYqgE4LeBwDj4EWOg
Qam2GQ6TLnZKgMJEF3CIm9cl2iqDp0XzWr6MA0FskpThI3pFN8e8l70ji9BorpXf
eqM9o8cJ8J+3qZFjoDQ7TyQ2x98RLWARCB5/IMN5+TJbsFHQ27EKrgIvxaFXNIG+
wscT6odA716A4VEBSyuydEMeBvlXcShE9s4MSReeeJ6UklNyQROI+xwNbCTfX8VF
bKeglHtUKwdd+VzVrHZM2tEV6CXqxySaMJIP+qWNrB76qG2GxJULKwmZN9SEVCOK
Dsw3mcw0Kq5Vm5BZFMM/cdIGBsxowooaheV6gUnDYsEQOVQ3NwQwHOAq+XFARbBA
eOM2rgUGGy47IaIMRltq24brQiNDEZ/tnv4vly6v0VXwV3+ANo21d8biEBkWjq0G
IFOFQCnpULodTYlyW++ZCdozSNUj+oR5HWQMHCQ0j7PN4L8u2Qo4gJT+8IbF74Wk
qetiyL6Vx0aeELHGdDkHhQttA5HmDU4HjgSXDhHvPmYGnCAKg4coptDMg4BYNQWa
GF8ssPrdNULPWbemlim4002FHpHP2Sb39mPc7TmPJBCiE0LpN+C/zCviL8NZQyBD
ALDhmQovyf9VVoEBCFUkpqDcyxCbjcvNtNtnZhbb2lKylk5VcLX2Pgps6AjiJ6wD
M2ruGJzH770K/MpFuvyl5jcwWfMTRUp26wPL2hIepmwr4/CDtEau1QU5KXkixsjY
PUgVOtcfmGpuUKZk88iAs7FNR1X93SkrOHzG5BzZDOS+5r9GYR/ZUzFi/7droFke
VWvtqe5xg2JdDS7rwp5mjyERJKb1qKo6tMtmfVlGoUVRLx1VCbafWIn9uQ2i34Ja
jUiMVqW/YvmXO7kxODNqIwCEN4MlG8pXNrwt+OwY3cncLFmL/jnQSaGtoXmRE8sn
Y5Y7cNLPg51vf/al7H1EvwcNxJ0SSW1r4oj4HO2eirN4iDI8bJk1hmzEcljU9CEs
pWRODiQh/YENKUwjIJuNCOr1Ngb24v7aGvAk+J5FGLP0aHC/qZfE8BdmDe8bmN6k
njeNf01+UL7sd4UVz5Dh68ojLzDrI4Ig8kbdm5VQiFDMILaIspFa3CzWEQtJLZNT
XOhhcnBcMzDE0hH9OCnqyCiO4mmxWwKusPg839By7E75Cr1c+UgmjR/3QIQ0g0yb
0VhdyV80Q1KCGMxbn7lQeKx2j3mtNPiG3Vo1VnS2TT8IyfAbnjy3TpS63loKU3eq
F12vjOwVE9Q3W+a3GkSxPYY2Z4MFAHGMpE0K230nulPXm4GU++LDINIZ3bWgzn5G
ZGkM4h85QvQja6TEGSxA6RhC0Iz7hsb6k275+D5w2+cjSPBFsrVkXS9U8fzR81GT
QlmjeRKkF5ARcEu3gEAbTGPTex7zsEOVR3XIEzESX9q2zz7O+7wuFQb3O9EVSh3v
HBOWjgcM8ug0Zi3nQRWeuOslL241vGbpeH40ZA51/PQofKL2VbbktjLBNqSkQQXt
AMQYcUxOTXc2Jdfe5PKRDQhcAPAehA52sedIZdPi1228tAugKcDW4O5mzuV7yKjh
207WTlGmpSL1Yl0Ja4o6osemDYqLGtXCSIbECsMc6Pweretce6kYcWOY8FcUf8LF
d5EC41vzLfhjpf67rukT9ykhcJhl01yoBEj7b8NhbWwM1kGjKAybZAjKqPuicfH1
VYKDdCej+awNe1kLzhD86U+OTnBxV5C6ufdLYEENgNxFtcUccyyqKvlmPhKkuWjO
vfEZORE7TNs9mGE6fBonWo1M7knRkQBF/ZKhfV0W7+/5FqgnLie/62d9rJAMEQoN
M3sPpjIMryi3cZB8d04plxGKjw5U3wflJ2sA8gMhXWCwrxZDUXqi1Ax1/FOxnbD0
Ho/9xgRseUPufipazZCLkMfB9qNy0YVfhDErbNz83vph3j+3Az9Qzbm6Amaf0NId
mLx/0j2U00MvHLr5hx64u8C2aUYDvv5zQ8HhHOVV3NMLSWCntlIljoc0eSaZ8jYw
aQcvPKAJpyVLqLu6hvzx4B+/6R6+5o/CQ/MaCuhpEneOKX0qMeRu6toxwx8KE2hW
XEjcYLKPKrtP1PmwWJIwSmiiOpDJnxai7TL/cM4YvVD5BSB/oy/Ma4SQK7htrKL5
kmSXvwn/4akgVdilfdhzVTGlxfETuss9irQwTjH/dxsg/jkt2I/SsAZN2aleqCwT
x74nHMaMNPz+9KlmiAHP0IRXb4MzExNlqoeLNGm5qkB9/WmFdWJZnp7zQyl/08MU
hXg97F/2J8GdB0UTMQxGREQQfafT3vJrNtiUPHCEfwJCRYCbJbLiEAU3HnrPziI0
d6YDvafC2sr92yexpjTgVXyPEFzbmomYih4XuxQhF06szXZdmY+XIMrD0v9w7MvX
YWGGMYa1yjtjiZl+63n7h1vKkxajdcjZ4CfodZmebwpj81pyuqYDWJKlZ2hDTbTY
NNQT6N/+8/pdzkOwcr8Xna1jr5htqwHF1uQOJkHRuf3IEK0wgwM3gGCtd9THRvT0
mrR6rZtZfrDE13CLsO/o9AHYDJvMuQ+C9pDnQksueT5nrWbBO1hxQeoJoaU+Jsg5
tm3BtBd4BO7At8pyXO2Dc8vxsPOFp8cbFdc64IEBtWvVyFn2XhfWj7kVi1U5oYd9
3ZhL8V2qryMxqxNmJ9j2JfOu71ENYsnox4AAH8OdDqX3wbQs1rLlYm2EVxvruI14
l//YaMwliyaXUt6/UxE/4iYjh4fiechD7P3ZyAcKdwqYqetaj52LMocZ5QJ/2yM9
jlrE9QdchAHlDKnmnRM9vPRIMsyUEzw6H5qlnQavQLu9bDPc6EW9HnWAFPl2lDDe
HcTQhtnkGjeUATe+QNxzmeVkpEYLVHqtD9C903TCZciAnoydLkz7mqLdGxYFww5A
C5E+eS0nuBLUafCFhjqu2PG7Nbc9b4hmrxVX10G5qN0/RSrGMOvHNs9Vv/0Gk5+c
d7wTiGCd16OXYwNDZ0oEtoAoLOlOuYy+EwpnAk7JGH1nMnVwNDfPKX88jGyy+Dgh
X4/3cwCLDRdo05lk75V0ZaOL3H/ujcS8LqLPsySlQJgilJ0Rv+fn4Bh2KGsDrRY0
Xe0fhICD0TnJKW0H35VfBj9sj/5xI8aKRjJgkh7KTD4ou3LH8muUSmIdO8iNgTrF
+J8nI7bUBLXkM1lJDJDHHXbaa5P62CwsKeaRVH1bdd9u9kBWl+AFUsoNP/E23+xB
op1QHK9/ue/IE/1fj+i6p8ZiDPzmywRm6K9l8U23cNC7LxjQhSQcQtQNTguf202w
TNrgUoZUNHO4j9FLEOHQlA0pEWNTusiYkrIUGN+NmJ/nHlF4UD/uo0lL2r+gdKtf
gNrD13c0xBp/pOf2ZrhDysiQYaU/XVtzeXwKrg58jefgBivEG3tD0UujxCON0oNi
aT0ZxkgXqqwGdYlcbL/hUk01SPLZO68jpUGDxm8bPzSug0b5ayfQJRSalc39Sp/z
BPiBBECRHPHM1DdMfxyP3szVJqIku6KsnJ6VyZNCkLhIpJiEZecNWiVj9sK32gnJ
GlsTXgwAs15Hqhxsad8s1Z0a/aexHQF5SS50MJXjzy3TGhd+CXABLvJa1AEhkaeZ
3usE/zbIl9fA82P3fg1/EEDvtJOX+SlRliysfORdc9GlBS62Y3KMpPDSvIabo5HS
7uzg+dnnMAmTXPUMPnr7uaJjQLqF5eJuO1uxOZ6SMKjA/N0LlwSOja9avlbBLrhV
UjmN92RErlpJN6YiZEUBxl9KVO9PqUmGQtETBCy+8uMHJQgMY9KzzIrESG7KH8WU
r6z45e53Hr6mVl4a9LqvzhVJ6t8eyUyzaHIWuiKroqv5hx0xB2iufDO30PLxm72J
WdZpd8UJ2l3AsU1THqPeXDbCtbc+8y+hgu7JZk3WgEBV8ok89aBdedcvvAGCH3U8
NMdQ/fzOI4XDDV7dAcuD6hTkt50K3TmoTmSyLnDw0xDR9zr0S2Ni0PUm4rOGfWUP
NPfGCdmwgGwsm6qLL8l9wstxI2k4HX8OoHXR6YdoEHWPOFvEKqIndMaX5swGblzC
tGdENIkMVx4teMlbzDHyiYGT7oAwJbuSbhZE03ZwHy/uUromm/L9Z5odt9aZ1k/7
lwI+SgFIBbfF4qV/4c6/lNMxv6Jlu/piz+W09S4Mfj3HK5Y1Aieh6QMHSOybKOGl
iHhZhpi5eQXwnjA+9L5JFjoT+jDwPcUVbFlSJg1Y48DlI33j1m99sdQnYHQCRCKL
5WrGyNtZHyGkhs1Bs9HjatlwdFY+3cVQblhsxtK2s+ENaH25Ii+SOpXzsvZOLWmm
rO+fDQj/w3cfnsJXxLnpAG+yk2jnfbSjRyf+BIb1MeiJOpWSKRVyQqwGz9m1XPKu
21n8cb0SIHcJF5QS+NTjxAWK33/qG5Ijnm9uFm1VRuRFCSuXjP3OCM8XL5mMpdz4
QX3epco0KQU6Gkxo+4Kbdc/To3cIzWpO/GUfkDm68Q0xgDJ1I5ipRwISaZguPcRL
SDQKmzo5Hk2L2W91x9QaGShP8Hb4IU/kL4sWAcoD1p/hFREy9EpF788MxuDYyGKD
53KsvM4xI5ZR45Sew7eAExfQF5s3tFu0BKmvK3ukjqSa+19zwj+PG+xFizrkiQkN
twljwJPDfJRTYLmkWRRYp0TSA082QboPxvlgMcvIResU/jaPxaWogFwMlJAJp/+j
pVh8aqC2dgFT6eA4rAKxG0aJ8ML2cRg7ZBhWQilGWCgLIc65AiIuisJYeTnOSo7k
o4o+Hmru6Gf9hXJtgaUR4o1p8ecZ3O2qzxDrkF0Ay+DwdsUWMztPN/KtptTdxdnp
TjPN0dvinKYbLt4aPmHVPSMwCwnebL5x9kqRG0I9sJNooKK6Y7ZccPv3k2PMrTK3
68obxLa51fjJWcI0uv2sR5Hy2TiOPn/H7Ks735u/OjJUh/Xv+90grHUbBN08jQeY
8J5gy6fykF63QogawMLrR943Ty9ffNL9XeGC6AlEIwTAtibqSRzgDlWgBSdsXa+M
Kvnx4mlEPx6UjQPBcy0vv6hf5K0X4iUt2FqWle/GPugZfUhhcwx/i8tOhuSKbdsh
Dfk3X7RzFGoMaypaTJ0u+isnCYq824oXwfWYt4DB+foZ3AcMyACYWzRUO+oRH+h6
lWrDShbuS92Iqy8xFReT0uEHV/0+GXjoMV7alfoahnihYoLVTOhDGYoemAAJ4197
7y2dPx5d0tqebNgQu2K3b/kXjZb08Ha4yHlmmJaDt16412OtdWjfiwmaU5aic7I2
cyMODd4tCkQCS5aO9PVMEFbCwKu9rcwyhQsEZ/bYsvgzufDEji+JpOOb1zZ5hBNC
ygFPgx0LL/fyGUE2sY0UfwwoMBHOG8/B/P+WlOhZItT0C+2GvciQ6HEvbOOb/h6P
Rg9JGcF0xsWZ64O0k6cHevNatFYvKX1F4w/mw97uo7a5hr29zKhidf8CU2fEchpZ
dKQSqzKeH2vGngTpuCnm+sMVs2tqUPvDc+yNmOu0NLnA8dQVza0BsEGPsjXbrZpN
Jf4BjNY8dVjXxoWTWxjvbGSr/TqTli/p1S98qZVu973aJTozdQ7crLJZxym97efT
c02jion7EdddmvWs7N1OgNylGbfyDW92CgBG9voIpRVUD9EUy4ZUPUNozxii+1YI
RHbvse2gSKGA5JNpixSEN1G+/wtuiy0o+DPKGx2tqbhk5al1KznX1IcKh9VGEuuw
EgvC3HDu+ok3JEXbyI8rmfSyfkOiJ6WM7SrmdMbbLaI7ag5QISMMAEkjvo/Ntz5W
tvDRCjpXQ3icatIWUFtWeb+CLUMerJhXBZPlTmDnO2mQ5OuXFhvxQEUN+M+4VgSc
+1frXBdvVC3QNBjxUKoic+5JPxqvMWnRt6qpkMjk9EPblqhT9o/X/wfqvtPUbJmo
AqHFgTIVS+cUo91YkpgrJSRXyVG6Md9+eJm+vaNchEvrV6ghmWLTHoMwSB7I+NHh
reyunbSqa9PEfHe+EtgZveQdSNqFia/3ZYqK2aTm9Xn3GR32qJM4yOm6ETuPLOI5
uIcFLzr4BR1HMOBPzz+PHwm+bNRmzbcqNNp1s9O8i8ODij57Y8SmOrPubPxZ0VmS
l/XlfuD7Bx/3b3nY1pY5OxY6Tbbx/whrhfHPfZM229t1PuyF8PlU9//EzxYmbEpU
JH/CYoYhyOXcYi6iDY4A6NIazmLgOxjjJLbpMcvwcLb3jQkV3P7qc5yWOEHPeiRb
jc9KbY04zmlZ7hF7mZBy8AOmrFPQ8d+jhPV7YGYjr1Z3GnJLTs8TXRJPA7R88VR4
BoN+uk7zG8gXjY8D95S/oieTjel2ohj1RUccdiVeILjBaiebD33vAV4b6hTKYjvN
5wYdZarGqEWIvKDqy4kGN1J2LN3NJ9fJf5DvsBeObGrzf0jFq0Txw5sROQzh35Gs
QpN144wxvBMpoeC/94S8x6Au+TIsGYvgcUTECWw98PSbzqGDyV3rwnDpuMwKRtZZ
Vw5JG0bCEk8WNrH8a96HZf2gMPSDsRBe9RCin4BHNVAuWrEzDVEVXF5fEPvwfgaI
caB3UQCimVsgZb0w4V/UwZ36wNVFT3DEX6Q5+sSE+DkaqCLYoeVlTjBEGdmdCR7P
A3mQKvUeytJPqv61MO0rr817wZFrIj4v+Lrl8VWZU/eT78H1iUwHKDI1DpZX/VWa
VC/WSHB8xo36gHAdqzp4Wr2ctbbDB6b5bxG8UbWptzHfsUZ6AyB5T9PBKeZOP7CG
jOxK7J65eZNJF8S00AlcUzKStQY56EU8RVF8Dz+aZmdGEM3gVF5MaUOGlVR7XD85
l7qXj5P3/yx/NTou+y+Oxc16sEfzF8ccKnb5AE4yWf8C64WGn8ytcd3tbrJG34B8
wnC+G5yINMd3jtrbxMGIRDAGgJinZEOruQXvtXU9oPkq17/uLqYo9UI2nn+crwY6
H7Sh5QDEZM9IcFe0740JnNSYSfe1T71AtX4vsQpQmzDb6LntIxDJch4Snc6GDwW3
xTHTzskPp8d8582Trr136XF/ZfAQbmcrZqbZ0HwlVB2Ap0Q1VwIjSULXZpe6dDE8
nfRbhHMec1LjJKpFvnWDDhDBXo8uH+zN4gkysNy+drDUx2Gfe4TQPK31ftneT/WC
NBOADUzaVXlxeqrpsqkYbaUwVYbn1H7AIID6mZUeoGcXGRRdwvFxMDATZVePSvKc
Li0GmONXZB8lMiaz9U+jasRmacXLD8JWG9dNJwFRXvm1YeTkW+6S8x17svrEfrUy
DcLa6txw90Dz78XwTQdtgxGt8bDSJs3KSQYulQIU9rHXDwcfJ3dKibxks80GjGx6
hUfk5oxqQ48ZOJgbNI9YjcshmWorerjz7fxtF3MVVFvs7TNHJyU9M7chypRw3EaN
6pgef+JYYFus+dj4B2q+Aj6+mZL/e5ZdWK0eV5UQsWFTGsq2abj33i+Te9M+AfWP
d2MBXb82TaGcjXfoDmW8SQ3ZLCNrdisTQIG5opCQ6W98ml7LYrYAD0B1r5wCpwYn
mCEionFRwT2SnW0kQ/K9xMHa/aRArpy+HUaIsFPSaRvNaq+sCHCvL8s0rER4M51O
en3ZWCOuWQihYxj/zQ1D9qXvbMs2ouMNN9guakqawAqooqAkOd+l88QxTdwhDSNp
YgcSl+wJpsHK7OxjTeNHjCia/34mlQINczplRO7KlOIUH4bJlsXbUAUXQ2p4eoOx
I/SAjoH8PyzR4ygKJUNdG4GDU5WJSEpBZH4Sw0iPzczwGTiLEGowzX6Uy+KCr2rr
iZgxlDBhqPRpX3klF293yoVasRAjVmDhaJU4GB8sTnyxBolSRf/dQ0fJ0bU+3gIR
GQFvCD/N1KMlH1vBnAUTADC2+59UKUPJ2CHP/1Jd0cGxpN9wLXril0nOOb55Huez
X0dA5lnes1hokivzUlyjTZQZZACPlUvv3zF2eHlmHGygiaN9Y3qRx05KGp+i3cQL
hBAcwaeOc2U1lWJ6CrXc/lU1rdoPR+e6otTPhi+6f+qg2Od/nck81dZbmIIGwUPe
KWIwuAV5+B7GSBL7jEQq0doA0WSz0vhmvJg5Ypv91JB4tGRQmHcsQcH0nDKCwPXm
mk5to+ljOEtQY0LGtDcfp+WkgswCnmr2XMGvU744+MZ3K5gWHr3ftYOQd5yGmj4n
/Z2vqT5GaPU+Nw9pzdSDv/fovOJX2hPfOZMEOFvo2yQdHtKk9WvSpisgDKRsUzyL
gDhggiXpnGf3Ikqo2Rj6U7WoehxQV/rT+pX0iB4Xly//0QPRFpKxrsFfy1mWYlJ9
0QOl12XOpnHhnNZQ87tideEFxXV2G4h0isUuxJbQD2ItQdXc7047QWIZRTr09Yqh
/Bt+j4wbxusWgXdOwwAOkwYeHpSyxtR/fd9oTbIpA5ALOFCCVkgBY8JDyrzhIK2A
kMTqJIdbaEHAVo91942mHFmcbFaRPUimT7zf4HktTNWFVsIg9w0h5Pz/T8bfPnVH
sbcegthEB0d0N1UD8eHFYsbe6vsr58GjKJYOuF6n0CuHYQww0te+W14vV2fpr3QK
s4bffmM4aAJNAJtGJkwPlVuYhkZR0WDg5CjsZstPDmH+tAV+p7wW7bt5KIS6jM2G
NBx6HwKOl/wOTD1q02mmWFd7P/wV61YZqCvujTCy21yqPWdgUoJQspAa/MiTpXPr
2sP6Yy8WL8m+bvz5Z7mxtjx8KMs/I4Es1f4AJBfIQBKHSUkWti/GcNUFuUyNd/dX
rVC/98re/aA4IBdKXEWNqQll8RNr3fp61o+suaR1zSAi+uoNMFHTTWwFhavTkSuw
4Wm9qupORKPEvEQhfxl9IB8H2kC/a+YPsf7aRzT35hXKVvEDrNxb6+nAlBqlhOGQ
5Hx1vRmRZKqawOcVxvrjtr0UVRqtVuhKgfiQPguCrBqanCl9w9a5a4SOGm+io/yb
u/YQL7ah45lJCEfSepvGxeuop7TlPiv+65Q1KBt2//psboGN7XoS6ouIUcCbbpdV
GvxjWqf+iGjbi23O07+BoE0C5TZNIzicVQ3DLzjWt1DJ6FRXuf5cfNJm8ck436fG
yAIavt8MkMLFI3groSaiW1MNKPZVQad9YwdUB3WTcsQpdmfqIzZ48srAnE20mFli
Rj29xlxBFQuvmG9xvEwGrzN+LBjrtrBsao1DN0t0k9m483kscRpQueoGbiDTcwnO
AkfUlNRKef2QIV8h8+ikzqeBZbkcj1NDnw11EWQTMxfwqxwxG5oqkCczm/cm3wjZ
Dvf2VbcKDMpbVRZGdzChtk3QD1mdo5AdtbCOspmDVUpLwu7OtSYn/nv09FRLlN6G
5Jz9fKfzlIbdg46zMXI7etcNUYmo7cS4ziCmtpo+gris5Cc4bSjFscfH5GIwBSyp
g31aDOxNUyWEJfCeOdtbVSL6Pr4EK9EEXeZz8VvpUloXrycozV3Ew6SsNjzP0+Ho
SJ4JprQLqM0xo5+RygS/RlFGIsszDCimW3NrLNvBB4TOHbV5PhLNot9A5REsm9xn
2U2cojq2xY0cy0W9zo0PxDN6JMIggldMs1i+JmtyNgXA0EuUUFZN02BlcbwPGktl
VmjW2jJJyJN4WU4ljyTEsB7ge67ht34fSDlmIWLXlGMMaKAJQtzTKAQCg4YqrI0k
h8vR4St/Vmb+RVJMrTt2dxk90f/D+ORjSR5A/x7BIdSSJcPc95F83Q8a4Z1uCrMU
jO1dCiPj6TYtZyS9cbmjUvUhIVY54u2OTgZ4+jZqGgoIc50ZiGejVkMxCT6Aqv1E
LQbpvXvDASCNrKjZZ7/2+TKYvSh56stWzsOs2YE0lJudH2X6I9wxx6TTpTGpwseq
TrL9N1xSKygW/oGvP7pSQ6B29Hrn4AfYX+xH1K+RzAcF34MZ5P3Kc6oGKvf27vXm
LCOBiqVg0QkRU2ll14PJofLIr2SoyV5yXwQYSnbrCTrjrqeAbZ5J62WZ6V91IbE7
RucMFeFNQVIiYH5xtrDtWTN2HJUicBnL86xqmqUd/vwHqwug6PBkWDr/4qaPeWMn
pxuO8RWe3vbhvQeAdlJdgqTwXCRerI+vGfGtIXHSolbU44gZI5j2xKcITp9p8ymu
Ai14Sai2/Is0leiNWjGXcO4ya65dXEW65wJFeie50gCiOyZJJddDmsLpwjhS2XDh
7rSZuIqxIdtxLeF0oAN8bYr96Sq7+vevDZpdY5a8GzPg+yn52q16wI4p6xG5qkBu
FVmB6LvdxbEE8XcVKKYxaGnBjVO6Xl45fv2xTWFdjzGLCFnsi3mEKqwveurESCWh
ldtgtTez5SdT9UB/gvHvn26si6JQHxdPMxkxOCN/snsaJQJ8wc1wFGRC6psWxfai
YFP7+XoBXbNB7A0hIhjnfZpxFF7vd3c6rZc5havhTrM0SbddDKjlCIX0ZDmTSUKK
bPlcph1Mmod9zvBDM4bsLHI1Suqk/S9+VnhaQXFmdmg3g9wz2Hyv4t5XuP1opK3l
5D5J+cnrGhzgg7uL+zM5GWiP/+zdoQhBaIDlRMZRv5WX34wmRhbDbUcT4rrElvdB
jbu71wC1D53N402Fo55zZn6Dw9tTUvFOhq/tF71fKvSCyu1lQubLf2JY14BLdV2S
bi+6PJDE0URxJDVm6vnzGJ//RIuvISSKiEWuAdkM1vEyuC15i8NawoMIW94ODsJs
O6cf7yHOVHwR0dmhZ9U45SVvupeUdHL5forFJDN/J/GUxfpSwonHEEulLwiyOe9i
OIkXZk2ZzJq6rjCXH2p5NYEjaY2wy6769K0xdqB6IbbGYAJ4k0K1rchc0fvVEg2J
tC/1lIl7V7DNpoRMjavnUQteJuuLk0pF7rXjebQjOXF2pldyyUPLNxiIYDkf6F2c
E1J/neUcFpXMStOcoezd8q8ICbdFXQrpO5DsMAcpedn/wU1X32McJBZOj8QEXAB/
AxvuFGMgFY07CQ8lefQ9E1YSiVwFvg7fOHF9o4yyXgh3eDlzhaz4BXgfVw8o/dRB
mGlZXirJm6thPazeEyUk+NPEIGQwaZVbbcFmJRRLBxDb0WywqN6z6ugqa3L8nXIr
NtWjCgAKzkdFoF0wuVjZtbOmOMQozPetmV5bX23YjNpCq1KLGaKvc1eU5RfXArs9
z38WD/phycCCQqU1esQ2JH6uidSwTn067rUKQOycgUSmlCgP6ZkC2LUI38JhRO3n
ieUHhjc+kClLBDI+2ZiJ//R2SlF5MLDHH0wNj/NHJikjlra+49Cidb1iI2ONp0/6
qYEIhLrFtAoaGSKkG+C+54NhXx6+USZQIZ+FLNR7xkobhEkjqAFK9z8sanbIlECu
hqXOALd6tg+DvGtIPudWV0rF/0va/KRnCScyT6OqmGxmOpSFIN/GUJQJlq/fns2q
woEWaWdmKhdwIWLpL8jkhd9KlJRyYwW53GZK0IC4IvAKsBWbBCMZ9p27XfqVXLMH
BVycu8bJkIaaOzIeiDEGfv490LkZsab9GUOWi+guMYq+lKMhMSBU089YnAR88pBg
+Gy+Twbn2kiI7wf4gGA5Tq46NYjpD8wcj9BKYcQAHuTDfgYCOtH+NStfd235fu90
YrsqVMzl8FyvYogzFGaiDkoIUl9aOAMwGOFsGl6cOK96lTBmpUz10HQKTxoNocNZ
phPDjlKUz/QCs+Fe+XUlv1Gnd3NgodkDmhcuV7IXNjlSr3ZMGzWczLqNEtbJTRlL
8CUlrExDCtRa31TQYVNCuSYqFYjJsrd9wfisOzwQZSVTY+RVV4qE1ot8XOL5CSYm
YvGnOrDIdYeAkJ0wHji73TfFmVMI7kavVDaOJJz/chSbW0EyoxGucC3Mvvyvouws
4jKcdrRrLivJw83VAqWGtyOzMG9tTH4H1mzpVM3yoXDRSBYt8Ne8OQM6Tnj993OW
TLMTCMAZ4MeAVQcz3p9up+FjOyIPWFSW5mToK99qhT4gnWTVSX5KUeFJwkyKlQR3
xHBkHGOVHJmDFbZbugGVO/mMASY9+y/+5vnqVrbPi8FvVgUcIMfbxEnali1FiK+r
aephZsSi4BkBSUMQw35Nsqv/7zyWy7dE4w/uIWBLm/zV4E4uQaXXKYF91NgtmBXJ
NqYHNVB+XQ/xKD1IGOoWRPxiVt6Dp3+oz9YchONBmAvH2LrZEohK7/p6fVQLE2Un
gGngwX0XE4v7VftLJQd15wxlFpz5Vq6R5u7KZPLnLyhfGZzHxLYTXgtLx5kSf8wt
5UQn4GrtqCaH5ilJ4rRvH/EynMyl65ym67DBvoPsrguwkIAfe5aRbz4+LIcOUuEC
2lopBc2VjgAJIkPv8TYhFxkj63HxCH+T6YBrKbm1yPcooR/5XI1qAbpP1PV+n5FK
kZJU1F7JH4zU1cygN7N61PIVRbeLMkqgYvDPTeQbiHM1Z6uXDzthKiEtlHECoHqt
vpdtgVn6JUpBde9lkF9N1HTIFw2rvVuTjbkRgyf5VLaNhZ9NGOaeL/UDr/0CZ6pq
eJ0I/q60ywz9vbOcy4H/twRnyrxNqk7aQo+iXdRDWBuy1T/7+iwJv8RRUPtm/H1T
2JewP01XPBvcmH7bZ3/0rjaCzbSuSZuUjuesICaxKAvSGPAdDUH+4YGeOiSUCK2t
ftGMJZsSiioRAAx0MnoNzd74v0aiigZc1+coKhYUK4aM77QywrQNJemniarM6Q4/
vWRtFhSiPTVfAAahCbmfeRPAOjBDKb+sMnmYL2CMnrB7XPoeHPPTxSeF8EAQczAY
Kd7xcn7WvlwAi3ocUShlWAOywRGltvs3r0FXhRYD8pS7zXpkTc8JbSxiSxnVetBZ
Z2LJeY1lCHqlSD2PgjZbFv7ftNWBqg2RK2x27RHh7qGSvf5oKxJVJT0uv7iNr19Y
s8TJ/L9DNvk0htQ1eUdyzesXVgdbBy4XPL1IxcU7bI4mPeGMcTtNAGApGcPlE5sP
zAtziOg+qeeX8I0kaRMRaxNTeCg5B3EPM5C8w3dG/j9GjTgUNld9relkTmhHU3Uz
U7whsR6MBor6GFwrx6ceicvXruzbW9ziQQqkmCM2SLxPi1NswtdGDc3rRHBxy7O6
vwkh5euNNYEjge+nXvKAaWOZYcEuD1dBEsE+2fq6mmDOOi+kO0VE/0d2lDqVFzgh
kAaLVJQCvYGB1QIbB9mA7A82TINRoBmbv9L18UEKC2ZtgvVwUY0IaL3z5c92KGgt
T0YphzG2KQbP4JHB+TURPhgtQyaPmWL2jz44tngY9RYWeB5IiSABNHPJGEE5HYkg
wN/Z80GwgfN0/YB17a4fqQnwKXxTqg9A6RzD2dXf87ybil7T3tjBXPQ1TphiC7eq
yeEAcVimDmWx2rW9O0xV36XUovR+YqufP4rlzlM97e6u2TUzDTcRaRho5rnoL0Q0
y69HUDvgFGirNGycj6sTUMHDNqxl4mzKGsGf+I6YPnZioZwpvwPTh7skAn6o8z2A
FOGQ7bk82HyZy8QsMeWR7caEywjm16C/hxa2qaJMtLHEEBLFZu32KBQY+bwkcHY7
TLta92ivqhjh+sle6vSmRMIp5bPdEwHkX7GjBHL6rIY1kmwH1RJ6xkuBZqNUSQgi
Tcnq0aEbusbH5AtmriIUzuJ6QmZfH9YbSouk4sPxLTjXvl81nyvaSGakNsC8gvPw
2HKO4yR/a8tzS15Wv0lduPk+QP49Rt+H91JO3fI1vFzJ4N4ObAJ2uaRJt3AkiGGO
hEhMhQpIHHOPShuSw1h0DodWZXDcVMNAaG08TGcEM2FMQdjemPLIQ0pcF+76eVh7
3Kwv+942NOMw9TelogI2V+PPOauz+dxVEq1/vWHol9viLaldxbpeYIY0oNACYs3T
oXiiqKEALRFl+vQ2j6AB7XYQLg2A4xFWnkkHgdHQs6XtA1nhGQKrpKrMtcxFSamR
k2QdljFdG8UOABk68cyHsPo366nhpHXalj7j6M5AhAbQbjKSfjtg9eMNGRLBOIT2
65hT3WNoHZcnStJvLxxEXwS2Pys4p8s+EzZyxyw4TxMpD4Yoqe3UMSEHiViDTlPs
eaoZSiExg3OspYRjH98YpLkVGqvIykGvcR2RQoq0ulFLHTc1gFOzt1VNGnANEF7F
MorpsUngFjeNTRUP6Hpxj+o0a9f8sh8XLcezIup9sw/Rn3zIsFRZyNML8XsRy5YN
2qOuPmS0aLqWeQ/j7eFDh3m+XGcs35SWqrmvUh/+lsSplSfWvnMYIhAqLh8IN4R9
pX5l7A+QNYzUTYhGqlGBOnI7fk4FRk55lXU/FcrV7q0zmFzM/UaszTwvQiGPTdRV
ju7cdCzhcfv7A03pPG+6cKzFuVPKfkYF0avnAoqz8DuLtZ5GMkpoyM0cWudWlSzE
p76eZyCRuZPIBHj6GEQkFbvQQq8I00ZTZ8TpmGl1WoxbCL971aP1V5FwNWi9zUOq
ObhN2FRZXuxwfDF36c/TEASPp7K3A5KExUu2/X/jvb8iignVtQGQkHL1JcI2D+uR
P+5D6ECNNNocfeJA4BOs5yDYLTwQPTaUvFn7tjT5Lkeg2cToJNL+KqhdVXqW5uc5
wFb4Dq0/cqdXFLfWQvgBerUt5YPl2NgNLVOjlFwcC70uQ1MlIZbeeOhW5pjK9q91
0O1w0cBXMdrupWlgxvtPFrq+IcQ3Xo3ywXkPnQM3Em2+AOkPis6Br6rktP/SmOXo
KWb07uW1Qmxwks8QgfXjpKf/ZO2gv9A9L0sMAjnusKLxFPaSkULMpbNcb0zCOZMY
B/ewT5K6Pvh/I8lJEUsS7Ah6aEePmWLx+vDZwE9jRjBsqgZBlRBhetJZCOwVJ3vq
Lde1v/HYtfqQVnHdsfVXjSPU0UI93B1RI+n1rs7PZAVmTo7JVJ8ijsvlRT4AiEAf
gBtq/1UROdkSb33W3riiGtgX98CTunHZdW1mAp6ySnR/HjNkToW4EGOlNf5C91Wq
lTBtUOXe2QhpnL82cav7N9fgwthc6dhlIls38eWuZE0v2bsffTyPkH7gOY2Bkvs+
l9bl2pM/BsqGtSAyiwye8AWOxQZN0G8z/QOPYbB81M/wPaGb40XSeOVXJlM4okCo
V8Gkuwq/3OxNH3WugPxUmaTXp6k8fEg2lnxcGGIQxfbxhoumFm2nWqCkXF18n9yP
9+hjuVYOCP8CnGiRJX3m+jUZjlgO6h0q4rg2J1v3O581QX1uF0rPseac5sX2vY8W
bTqvu6DptPXtxRBQVtUxAakP80SYXaJDkfaqpA3Dv94AVoxYKDxY5Mj+eFRL6vgs
KwCCPkNsED/HA/KekCw0DhN/l9AHwhdXmJ561zodoVdiqfFr4GRJSRD8z/9vBPBE
67rtK4mlddPb8Ru4hp1ZBtz2RfAf5JVV8jEZ9xG8pgmQZwNz+vQnSHIGpm8Ses2q
EBHHJrOWqe52vHZejuI9dS/OxzvreI/RJzOGDaJ1nEU+m+OyY9nmYQa9iREOP5pW
JvB/Gm2rj1mdKz7TACuq22mDKrN5u9aRrjVHthWlpb6oRlGKe8Kt8AZ89QvgFqzl
EPLDLMD1Tsu3oO8O2gUj6BWOMjDjh5n0arJG15eO/GDXYG26j5RaO2YJvqqb3iKy
AEWxDkZ3I/9/jM2WxbVyaRuVgcT3r5J84IzGbAEgIcJttKrS+522nwqI1v6caFXK
JyfiINcQr1rRiPOJx7241RZO+/xiaUsgcSeL67XsyyiWSKP0mMxgRj+kOhKo+ycC
/fuVVtInRSjYvXXgxZdinnAQC/4N3YFh6C5/Mi/I9ggB8qTOhLlX+3g+MB3jtSeg
eDZKSwgVChbe4j8xHHOjIbl/0/B5HOnzyFTktU7Go1aQnuZSlL6t4JVVQ3AGtJzr
ql9HgBe/k4RXqbNKqwtAdetn6acDgWXt678rZas9zJKem5gdazfllW+NP04RGaRR
Nc48/V6PmCE/aPP3ZYq8j4Br0vFhWjswPUlYWeIPf2Zgu4FUf/zv9+m0gsGYU2pO
occsWLFMnr//9qMt5huEI64GsgGZL6FikbwyMk1tFHMm2tI8SmMNjfPULoxxBzKH
wyycDs70GBOzC0zAIB/XXZoqxxvC3Q/4uvN8cvEEYxb1IJEeMEugiQgeub7ALmIt
HS0ds6UjY/n/DE3r4O2cCKYqyacenHCwJFLy0TmAT4EWOql0RbJ4a+kKj6eMTkff
gSLQJIORmP60tYOmNl9ZCIn6HnkzqrGwV8ftuvMl3tcRrJHr6jhNjgkOKf6XX4vZ
+9xhpCyJSHqKiWjctd35CYl5xHOlOcIAH9P6y/nngcIjFozpjYllhXwAJ9lSFW2H
/T07Jds24j8AOlbqKBBUz3Hdl0h0lQxzIFSP9T/tnAT0Zshk9hF54SQTV7F9cjdq
ja4Ybm589zvn1XJQ/hE+ZaOcdDiynDdnamjb5FPbINuiwvV0+s2reb7J35t8eMYd
pnO/gCUzb/ndZslr95o//rVczam9MYbW2GmD5VPuj+xxhVhqRl1zGFzgv2MdPfLA
0d7YCUupoCW9T++vKPpisP1+4zhENX/jOOJUucPFE8NqNAcZX39n0IS8gNnfSpHB
JmfbTR45XuRqFe2QRZXhEMP0GV1eubBa3fHXAmjZf/uGtWNOLcHXA77UChGZ4T8q
gEZ4gqcbf4vM54d6nT/YUP1eSWAzE707B0V7g/9O8EgbgUe+zI3L6fjA2JoYGuaL
D/ouBKNZGW8/emxtoqjPlLefylaqZC9va/0XB80be8XPgZxmQjxcYJeFeRl9ptdV
uVMWbK7b83Xoi+cV0Mahv8ryTKTg64zMlwRSOdSCBhq7mf4AHM1nkc2EwCxbIpyp
J00XgdYmouC14wUJ9/pWC2JZs4XNFg/sHhR2mmepBMSZhYhcdAjRLxnaN37Ge5xB
r9MHur3RK7a6xByOMTY5ckZyiUkp8b1oA4BHpeIYVf/H+w3ShuXJDes/jJ+L83FV
HowKFheVez+/nDUYQ3l8cNkX1Xqi3RajGUZChE/iJ0ABvGjGwfy/PCZP9mlP2YVu
rRDvW0aSNiGzrRnf2/6/FWwoPyzEW150+/+FtHPIQgFHHYGKq8j1COJgF6eo7xTL
yewTdjUffu/Q9YpMrSR9BVyZolyurbqOrrPFSFgQcgYD92MKs7PNMyVglyy/VipI
mVAJA5R78IyYoHrNuX4EuHOAgiOwOfkj3zVEd082yyUwMmAKxIGNOg5i7g9zyALx
4nf1r4yXjWAn2ik9FO8S74/ppa04M5EeScsFAqAnC8CAkPl84WSvd7NXYmOKmW6V
HS4U0tKoVsoTs/4LQZ1VFZ/cOKQ1iphWTn5iMELjVmcX0qQ42rkMy4x4bwcPWG8r
r/fA3z+LOoqmBYUxp4YJpfkySa5P6OhOX5VOZRMokw3vOsXCoKwKR4Qq2E2BX0fD
sJP05uJZYmWalCdEdJ5zDDGqXgjxUoLE0IbuP2bkZXlGZ3xLTlsPlt09gsJJgT4+
UDvLBufQO6B0pdGaQAvUOyNJI3oDw3tU1QIDkJrJe/j+pGidmoFYkIvU/RwyHHrX
kSpr13cUyBSgflVVTmhDZKIAgSy9M8tdV7ZuPyVlEbFabpFhoaNG+EnVsNPkl6Xl
1FZwNab4qCkz9Idcj/mWCdleGq20S5xVtesBFq2cPfXtrGLY7Qc0jwbdv6jAs2wC
l1EPF7ovKfVLQkkK5rrPwZv4hYkDQj6gJwruEICKpiALNjQAtegMLM0blqQpXD65
00unWhjejbu5HvFl/h4UyzghNElHlJnTxndG8vbt/yYXXO+T1sbyNzK/ca7mPvl8
LuHT0jJHL97D6WR/GHqIwQbYbGFOibgRJSJmbiFs7Kznv160cdEn7RYhLX09OUrB
GSq0ZzOY04onesYCgVBmQGLFGFtWsgqMzJrds8aQk+KkisNhkE6ahsE+CiuPBPeB
cGluaSh12w3LpAHiigj60QINZUkYxulCDlWEWisZZaiqxRseIHFje6Do1HtaWqmn
oRiGH9l0/6TGS+aB69fLI3BCd0DOmtNYSY0TiYgugWGHUz+1oJEamXTxXCkVP0St
X94Eqv+x7O/3PPnUV6J7QnstdXFPIss+YYLsTpsaQ7fV3uYaO+1d1LOLd/G9U+/+
ES69nItZ7c8no0RofFP522geIrr6Zf4Reg7+8arcleiBMnr028zsp6Rz6whWa5pJ
WFW6MfDGnXmT4lLfjQe9/4DTK/wyNyr3umGklDWWJfaC5pGvwU0tnMC6Ac37gTXB
vaqAwPgO8vXYPvcp0trI9CE3QRY5IvGhpuhEC6vPxzm0AyTJG/0yQ3EVlT84B9yp
eVcqCGFoRYV8ygvO4ESL1uXxRDHOEu5graptUGRE0BfaZwvgfdXxUD8EpLudWScg
mfC9ceR/HtJd4z7aFNmat2VFLkW19nFAr36H8aT7ZrotUQ1PTnJWKvOBJpUUgI9/
rJ+MQeDTRYP9rHbg49aAg1KhMZgMJ8xLOwc56Uz3vGLEmgaiQN0JECZNq0cQ2gLb
B4uqNGeVmhvOBXyyFl2OtKekCgCOKH+xl8UwjbbwVGKRXP1zKouSXM1vRpQei6fB
A9WpvEi3qAyzSJT0YvRJa7JhglcQzFg/wmrBNMZLAGkuwgq1Y1uW9eFu+6vmNJaj
D20id2xRZ+j2oMm9wWGqWpzXSXCzkhRmCV1HFs5hxM3t1OHnFMoE7r2KzW5R1Lim
52VPnxOjJ1zKERqDqzIsJQWRJvo7fyVF4RI9O1DWXcPVHs3Oo8Gm7el6wbZaKIiV
9LoIIa26LaIljmArLtM1UHBMCL2sgUkERftUhwmHpSD2w9nyQlPfu92fJMTIwd5E
9PZRAT4HY2nZL9ERVqAQsk1cgs/v+CqoVc4L47TGVU0aCePaBs5tIpfJoxnoDtMh
frVwhmlzcrTPFAUX9laqFn6RGRKGbundjCk+Q6eBAhwjQoegCMWiktCBnfTA3ddV
U4sg0UbOwUoN4nfbsmMEXA3yZze60ueZv7MJkx/iW7uv72EwQ043P52zpjlhcFCs
aiaORjHwKJeOuIn771xpdx/5BPVZGemmXPCqQjCRB7My9vSeWZbLMiIhFntAfdAk
6Z+lg01SJpWTI2/fySfyiJKm5nNUd4L7i+bxvTIyzxpbnOwg6ZPjCkDg5pT84H8N
6jCAUTzVEbVjnlkDOr479Ir+SdB2fIa9TsBZ77d5Sb/Yat1JAJQ0vnNvTrKqXCtX
wl6/GVrQ7gl7fWhyYFEEsxGH71ez0swt5S6gOr4rKCs5oluFTv1zJYXMD2eNmZCE
kLWMq+5kKii2PzPbnQJxU3zw+NjehoEF1XZKx8v6EmDjXnV8S25XXWyMdyCm2+14
9wuwpLeFrGtw4UtR2xaRogMZo4puVodkFbaQFg1h9+L3LCVhVal9TX9OJHTLsZo4
pADlXuLf8nC9XEYAxS4oVBBylGU5qsZhvhCltN3SbklV9Wn3jvXOKIE3UWgqM1zi
7V+iZbpI7eHYPu5DkXRrVEsOi9pegVUvoTitI4WlMYoH1xs+AnDzo557SrygOiQV
Y/AVgm+yvtkr6scx4MyEZfxZ1E7pwU6mpcNglhYr1u399I7iNqfTjdCNMGhrbrWR
z3Iha44NOkRanbp+GfTzc6YiNzmHApNmEqSBBelsOLXpXgFWVe7eE1KrD6opEvsA
afzu/jVPfq95PzorR5Jjnms1/uH5R4qWVzunL3//MG4df3Smect2Qndw785VAUY1
JUdAvGDM0N+IbdnJQgSVcZKm5z6Mm4XGi/JVwZiXENfraSMOkGzDt0oDb8AeOU9J
UeaYJ1Ig6ARAv3Vf6XmRBPaH5kKfnLKc3r4iPGuPO2bThk6jqnUQ3jzWU+HBJwIi
mjUyV09lNoadSncZdw9uxoZ1tt2xP1H+R+7gyKbfMOpNpO4VGI/bmMRsYgcjz2iU
PEL6AmlHOtKNOb5w0qna9YieoxiSUJLpNvEeCls/evuNvk4CsEcmN4GYnUc8T8Qo
AtkczpymHOHT+tuk8XFlrWhqqUYj23r+s9RM1YuznRT1a5Z6VwO0dLi8fpa3RN/4
Brdg+6A4G8UhCSO27LF9QRhH61J4NCiejDmmpXRZoUcAaBGwPgeUUNrxwwpQ3ttF
m7uQJ3bWwjJd+hWdl9FYqZxPEmoVBCsKOy8IVg8sQY0kH7pVyqpv598DuNcsip+c
8Wq54DSwiOgoZPzOUiQO6fng/+Od5OEEuFBPge3BpzQ5xox0WTcKZ1i/JUI8YcJ6
dKYQnZhLVjmxsMU3vi7PMXw2OxlEDKIIQOOILqSHvH2lcy2+3igP/cFf4zsfv95k
mj22JWYdPJGsr+JWg8uliaPsgxiEp6Nz9Wp9afCrQoSXppVnU6m4xal8PWmWruuM
yo7huf/6n1dqj+Z+IDmR8nnpW7Wj7LF+Kv4hI0HgTKv32j2+xyzBhIPQBxrbD57S
L62Ygo1P2ykrojXQgO+FTlY5DKwAjQwJcgLwrvHo5UmoDwhBDyshCiQ07gpjggfm
T382fB9ap4SeJfWntvnPQ7OXCGxAEFDWcr9LwKHLSZpmtVx1iHLTz+Wu3MEpW9wT
SqJ44PlNYC6uz3KbLsHJwqQtFa98ZBoADo/CHCesK2dg27FiARp941J9lQO8WNiV
BR69CnvEx9bPuoaTBHOtu/QH6VFqFmzyp53+Q54QtrbFjQhk80gDH9an9nBzhhXE
nHdpdw68ztcKiSP51oveQZpdOeybECGG/gAjg4Xvfy3z7gYWwN8PkFA4VboglhWO
CbOISngG8Mt256NyZ/eedo42AO8Xc6gd/fSD5GtculUDC7tHH/HDfFiUlIRSMAKC
A9qkpnpidmaKD22kKPCxKPWII6tQEogpg9PN5scKFq2BZxQO9gBWf9aAA7gIEzMN
NsA22qt6uym8R9tX/d25H6TkUawbliXCt2LnAiSBrBjIgSc1e0v9roh+v5hIY+ov
CqqgLbetm3gIEWfsCfeDLTZ46BpKwdifLvEpdcPn8nmWQz6YfkT8fRZRPkYQaGlw
meaBuWp9RN0BwI7ig/SDm+eFDqSLQBo5mcn3qH3ViATqFR2tb5130gHZvt324GKG
TayTOx5xc9BaIjeMJSKYaII4zYSMLRjtPMQDrW8dCqVtwNUTdhwFw1cN0t2TBuX/
xpqGCJzg5G2I12cqEDOL8/rDjgKdarPueOqXja+BWVsPmdZS36fvSEAufJbMaJjY
pP/OE1IVkb63NaV5LGnhN92NLgQtN6PWJGb0vEMTQtoj99TnDcpDaKsOZd1207oX
AmB0kwDT506tqhFwrgvUSqJCaboLcoJBPD4RWWqcUcHQaXpBiB2aVpM/CeMHIjca
7y5Nz6xJVf0lcdTX/U3ifnq6D+JcmsF/oWkBYBHBqD7Ft32wjBn3knDU6ocldtnf
WfJfLj6nx4f2YkPdPIhLw+5kQv7rxMy/FeTfy7DH82MclWZLKvV+HS3KbTJ4bx5X
poKtRk4p6Sf3yGbKU/UOjVNxyaIHvVqcazQ45odjD7NmPcpUu3LcYnxEvGX8MdDq
dO5BUdd+UHewxxUMD7dNnn16uCTT2ghhJMHK3brbdp2O/g6JEcMhuIOaYQPDpzFO
af6im1Vjit+egyjxkcocrijjB/PiT/MJebLhHXaAdGLEBWshNUQN4pYYByDl2Hu6
4iZDVjrvOKgDnxyA90qvOQrYZQC0crtG4E5v/Flzyk3FFuJrwTsVyIqG1cAHjioZ
zGi+FKQaxphgY7q1nS+WJS1BzSdnlGnVDUflKblqewMxWrNyc7M7jekeIebXhJjc
6pFxFNhLGh/Y7YPouochJNbt45DDqxa54ivwAe1zpR7PdLShGf/0iqAcyhM2ah/9
zKs3xnqSvVf4IT/fu6uh+fJpLwVU5xQycE4M9/ZGaxg7IBaVysDRo+uZsgZkWyQI
cjFCCFwOS4r/uZt1nfzqMmHw0pafIkdVkXHGzG5hSRWX9XlpmfPFgkm02eMBEw1M
b5jiBQYdtczjVxhbQ7ddJUjiypQ+i/4RlMh6SelJ0zCMica9UKqNfz1RODv/b/AA
oIpg+Ll4sFGtW5LeIKQtD/vOofJRyAWi0Mw1CfQr7j5dOMxkfbKzA5Zk+ipmulKU
YNVPMx9RQjY05n+VzDTU6juVJnEFOzHt6wYdfj21VNRcvafZmTa9I2XYVvBodcP3
aj2zaHOr0ltgj3qdqaPmeHJW4EN5Vp3bxvC02wh0C5Zbbwj3wctcbSVNp0d4ksQ/
uEMWxq5PVnnqgXid1u2McdavK/gsl6o+i9RmH817XlEYRiIn3LXPk5H9A5vx3l1y
8AWtcklQt3QYexGw17QwywjGedT6GLg+noYaj+mM6ZfqduROm7odNxRAe427RU8f
HtAIrHMJkj1yI/NuCgVC/xdK393r0BDLem/oXLO6eVPsz57ZyMRxNVBygPMZ4tpU
7KA/z7yfBuUGTzL99Ssp3TnBa2XDB1ZrtxQrCv9fgkzONKNGSMdeQuAmbmA6IREC
BWccsxYgzDZNgxoW5ZDRIAW1Mp24eoqkSnVbr0gyeyFsJdqBmyNlyyfSRmpBi1A7
bm50SAVk+ljXc9KXNfbWAaxlqBc+ym7gbAnI/mRjDpTow2x0+JqHQO5Wd/jlP1eI
8XWHuatgWK9WwUnMoLdhv5TVBnyCO2obCl4qT4zf6lBTI72l78rSB4p502SVUhko
BaGOfB6aOGwQOXJv4XUkgDEUtG+ZIiGHUKHqSvmP5ue9T+8ZDpvetgKO23bLydxz
MAI6/Fb4nvenbxO3EX50jlo5q6QQ4614EMUz0NOKxZnnHilUP2ekGETTANWxcOip
N/zobeBAn+4TgjCiCT8lHfNlcoGyVMXAJaQHWc+Wqg0iqB4HPB+5WIfMQox1T0XV
Bp8Osq/hPjh9llPG1TmsnnKCbX6sKq45iOzPEY2e9XSYc/Bs9nrXmiT5absLXYDS
Dd6yX9SZ7eEsZ8tyUUCMLrGGJN68xmHIjRw6YSAHLUINO15QDTT7DfKWcuZsDVbG
BTb2oy4ORvHWBTiKNIRu87XUF40hEz1O3U1iullq0rH+LD6B09E+xT8Xz7dW/NeO
9ndhRdF/hUZwfp6lGqtEuPeSzIXj3h/2ySWn+RfyCsYy33WNF+shmcjzbBFKcHZG
LSo8SehjQcx8peNTRgJTmFXg29odJezTGkTWxUs91oxBfsjKVP/WZNxGQfKY3U08
LuZ+GFXhZC174PFBI+0PpZVn/8HGxOw3nQmvvr4LnXcf61BJCTEkZQswe0PykriG
0TKXk52KRRpZGcdIW9wFt1JQ19kDnsjEfKz4PCKp/Yekw+Fxxdy+TKixsc/hZ5Qb
ST+d0kx+QtLoVQQxU0i1Ig4LCTHs8Rj+0ux1cnk4206f/hlWgDfRdbkumqcDoPpd
8ryoUn8u43aZWa/nuu0Qtz5q6eUIMnN2SJT7EqzUXBwnt16ew4ULWyz+zKJpD+7T
XIUYRg6phw01iUeMA/3CMDNsl2Ac2DwXledDb0kYO3aI/SLS1aJl9RaYjciw37CH
OyELDLTA0o0Mki8zVot4JW8if0bxqjMmfKNVZUl3q1UYwlKA25py91E1VQL4z2mv
C1WKnjjheJ8aoirkU3T3NgutjdwkNuekaWP5Ozt7FtsntFn38rVC5dYLoev1StbR
3PxLoCkPJsoy6GmHFitJMtqB7GEyviU/dF0kpG+Wgs2tgr4uxIz+5p9XAhX6P2AF
X6vISEtAlTB6BVWVt9udqpfOjfiAQ46d3U2hiQY6jUtyumbOJX5k4ZGFCAxz0Fix
vJSW3zXihBAJbAl9DRaslwYAO4SYVUQr3LSjC727LpmQ2buP6B88MCv33rmXFT4+
G+8fSK0YiE+8wVRRs5cNtXbQMU3UKYwuHo3uHqzYf1JzwyyehJhhTeFBG9YYJdml
25nNpTibR4lU0fbznh68itM/r5qF8g+krPTksuH2xn5oWZureCG8EUsZ2yTTtsMl
sUDM3L3DrTcCPWdXBwiKE6lxB88usRVOJewfSreovQkVGyYKTh61D1MgMmgcIWNq
ekqvY0LBQoqCXiIzaH6h3rriZxSR5eezSLg1DSqZcw08KO8j89QeEDbblL2JdBvd
WO63xRDdcLBP/51lCX+clYZlgqdBFQ/tPa12WmcacY0L0uB8CuldHEH1z8y4JxtE
eleev0Nc9X3CXo+wZyUNd/WcYrrG4fL4BTFBv6s4uTky9hlaSU1VtQktLDJ4/dsz
zO8PZGh+oynOuy8PlDS49VHX7fdHIdVmfshjWMLdhhOqHT0aNkljyJNo4wBZj7VH
AH3lTn0RYRGyKZKnMFHb23eS6fiMw3nmQ14bVeDYni1cc908DmWdZ29lzzxu8+g5
LcZTn9K60tXo2SX0d/ZR5C/tkIqTQFUI71FdfUviqqggn0JKNRV0uxJVh6seMV6t
JVXHO4ZwkMcC+WSdEM889BjaK5oKDTqxoB+N+Szu0OEvDXV378sUyJw7H0CVOLeP
XVG5ooJtOx5Ird5DuwK08TQSr2Of/VlR5kstBq4sEVPHspaiwlYI27IGQDJlv9Ah
/Mb/X6T7M/oHwcBV29yBulSgj3JUVjpIf9rGi6M7w+laCUGL8lf8tUXvKOWncxlv
xDrAj5oyoBazV8Tpbi0BzCIvJXUTwFiG3713YwySkYprnZz0CQwZeGwyHYvib1j/
ifbfPuEVZLRQ3E5FjFeHXowCj+QT3Qc7f1Of9vVbRoMP2WGKZrdk1P08YvsAE3g7
BztR+L8ZkKeZ0uhcxMDyGYy7+WZkK8H4c2KPJSwvK6d2kj9V6YmntCMS1RPDgZYA
6Muk667Reil6EHmVtRBgvQYDLed+VBijUK8JhohP+csbNRNUDMaRSCDE4LILUryq
DwZRLMr6peQRzLA9o42JgSZNOXNMiOAXuK9gqi6NhOkIegvZb8PrGtIholrM5yvw
RKemk4TBy6ugDGLcEi3/79g5GIPqoLjUgAjHI2tUyy/Rdv5jRLCzjdC0Kt8H2Yd/
cW8bPwyYDqAEeghTAn9P1amsn6Hxe27jt2l6D+V36umHvxvB4uu87QnGDAsQ9WeG
R/loUOlauo14PArE6KtupB9LjY6gnn+aTsWjUdUmBnRVTaRHGjDm+qMjRsWSHv3A
2spkD7Gd9EGIr1hDWw/ET2eIaBHH4wrYpYyVgGPoBPvLj/+2c2MHJkcipOUP3dJA
hw8ktuMeWx8y2LD88MeClFwK5GvqNxgfDqLn1m8BXwpbBC68qoUEJMELxwtpbESr
+QxX1ATfFQD9BEEAzCRPO/daV23clPIzzEHNDuYQQ+MZuJLjFIUYxrrPm1TSHKVW
NfyPagzmtk8pZmBQIetXEn9ghd2zCK2sgXu89SKE+L8kXsgh3MvRDfsmzoi+gU1P
2TsGUIiEuQpKOfSevLlgxceEAMZcEXhA2pASB7rHt2vAxZRiFRyM64/cqJCOe7HK
3rUiBPs/WQBA4XslJm4mk3i3zoy9oJr+b9BsmpM4X7n+gNCx8yxqltn4w3C18/9j
8vO+qzKXPUdHp6QQy1U8vAtUTALA8IJyls0WOVocXu4vk0eXpypYdYDTi7FXoR9F
6sGLaBg1oTvSzkkn4jw6RUSKkG/FcRZYNGn87jMW4WpdIMFZdR1Wl3OTbah6+Q3W
6KyMFGLOLvl+DWATyv929cYGIACZ+TgKQlNHxSTpfeAIilpVygqXT/EKIu2dhVEz
I5d+Beo/TuTPIwBdFJljKWywGyf/GtdZdTPQuac4glsf86/l8FiIcxk7buVDME5+
kyntQuD1K6jq9TOM+afvxnQkjts1fYaxmL/5kcVwk8PmKDxM0sorKWVBCVtvCg18
pckyGNb3/gX/LBY5PT5jYTBIMwtdyocb3yN/mU5u7SNMtGFu7vo44/Y2jvEmkU4B
Ez2i4ET7XjJG7kDNE44bUuLDWSocNrjMz1YYZg6mOM1caG3nVA2ahvlGQWbgNgp7
HQ1JbYcWHmrMqXAtsn8h0binqSqNcWvHQbn04WZUcvj4Bkb9JVACHFOQSMwooL0F
fvZ+nyn2sT/i6TLm7bBMfc6kEwpCIzFd2O4JDwxMQK2KKJ0INE1XoB7p55rGwb6f
xgCaEAMbexZidG9EIa1WpD39csEPCViZFZbn8XhChilYnu6wqEMk+Ok1nwHyGKBx
Djx3o7mr/z8by67WUYfjyxQ7u8QIUeBZosD3WoaocQD8qVVLUlN2pL2D//+SI705
5Aum3a5cq1iAjfMJdcf+RvAZa7H1hHaAsz4az/zF7sGGd5FQI3wGDzpaYn3cui86
GGeolxtkVvNFwFqMPIhyrfYPuDIA2enXlFpK9qbeNGl8U8hjjLF1F8jG5QziY5+R
OvcxcrzbFQO7zNpGvgcLwu6e04E1PdGvaX9TAk85/nOvCTiZvt30ZIVRehf7Os8x
sovNLqtU74VPYAEByN14wCEjDF4EwI/zUwwPi3RN3dacAFQo7V6vqVRPlE3eRz26
itUAKtGgPK4TdFUd1u055CyL9WV0CgP45+5YU71fBHrzwVJftWdyRO3Gp+PblZ2D
U0QRECTQf6Hy+p5pA661vaGT0FrZcMkElqxt6evvIBfZiw2bx3HpZMdg78as+H/6
aX6XjhADgR0gTfmS3ZFUm7ZUFd3QHpWIqnVsQ8sj6mO1s3COrHVKUllMmaat0zvX
AgOzyF+3DSLW430fN9+pSDk7Y7YpFSbpM/SQ+e2FCrUcNdqHTorWro4z/FeD4DOa
XHqAr5gvgZpAF6w5oQ/LcNBZLG5b/KXAYWi0lrMoIdfnK5YxMTbE+uxmC2bmDggc
zd3/f0II1/Wtr1T3zo2tatKrrJj5SaqfBUHkwdwAcjcKoJusHhhOTHA6yWg5U6RY
BzhGrDTloipmFE2Sn/sAXb/rXGavJ0TL/Zh/2LxBRU7sO/wdEfb9D/8f9SWisIss
3wlH1x+EGKwHh/Ga7H7btWm+vZM4VhCNCcS4sfapNitvnKpmvEtglFZ1Kb2VsVp6
S4xNPi74lY7tMMwpTJCSjKXGfIK3VbU9y3pLI3GL7J3yyIQrLnTPFHbHlfXcwHyw
61282ejLsuT/z1XzNuaTb5VAyfV+TrQR6pkE5rY5H63cWwSxuPJTuSrdRFpoyGBU
46iGgwhFPaG4o/kM22w0WzYvVvxWtBQiYmPuPnLADeGDgLz5aX310pBhIW+HYvtl
woo/tszEqLYj5L81bQKbcS/YqFQInVBIMuQ+HSKSZLoEpcs9itv1WcpcTe1PSloD
mKIzRRpcM3FxWe1+g6ui/qrVdC+TD0TgCPVqX7wN+h+lqlNSKw0yUDGyX4EXYFy6
H7vQattfX3O5HSSE5MgMl1mbwF72BJfp5Tl6VjizZ3GsFJ50KNgNS8H8rQVgNVWk
9nqnr9kUy2BONuluaY8+lcA9G8vFq7vU0Zb/zM3FOp/9ynENUJc2pa1Zebj6kmLr
IJhrGibPvJgUPutDr7wRJ6EZnvRMOnaeAU7Si+3OY/8eq3Txjwr0VMNVZvkux2Kx
euDfh+K7mm3rRrh4swljzjevmZPbpg1FdiQSjEdUnwrj69SnDbbT9SVKxeZ2Ebey
dXAMgauwPxq8yX9fEi0kA2U7xTDYlIA5ahScu6Ffhocl2pu5rs50yQKAjsynbPFq
bzPo6qrVf5ZYt9Ifi3/ioTMKxyEyg8RYL7ZkNlfFIRe4If3h53HtsooZ1uybdTp1
2zv4+QQq0GJC9wAAJ2lnqIksrMuTl6gIIySmHYfWyhOFfrcMut6HoSZ/LL2yC7XP
Msonw3d/zUvViQ0JOrlhY1Czx/d2s35pK4yeVvSwTxUqerft8LHyMGCE9R2RnlD0
lXD2TKdUZTLAZU1L+0mbk5A/W1qnBbKIQaraotC/jOL52WWL8xvzcIqhOFEB5ySH
LMZjIwQ3F/mtOxWvURwVc8t7IvJkGpxHvXoKDinUgkceZNJ709EWi/+JF9IiYOYi
WcRmqA93HEE1WSPvTvkQ6m7nMQYbpaoDzy8s9s+iDDho4Wkg3wTulnctjJY46S9/
AqM5USwvTe3dBKsIVWLDSPy9u1FwDFZfFgSsMJ86RPtCb4CeqCp5Tl63p2v62lhv
vF8wySGJigAVmY7DgsUvAmzd0DuMNu7gwtYYGjUKDoTlm6FbQqQrXza7G2oDr6Oo
RAZszXUMNpu0Tdo64HhhPtcLZlW3yW1xfzDRkPYjcSi2CRWLIsVkH4OKuDTGAtc6
Z7HyVeD5OzFvhBj2ePsHWTKn4b3bOW6DrPE9H+H6QQVKXTfG5X45Y7YbWmiunQOP
vLdbgMzYPyDtn+ho5j7py6rDY9bXwlC5GNYWruwcJWGy12MvUju2UE5lO11hAfmB
I13bACyKfrG0PGmc/WPXQifSt2vkD4KxvNSAEBtkfvL3TGMW74weF36yK8BBMa7y
CrJt2uWbaZKhUsvVcvdh6nF8a/nuOz9AQ6C0YCO7y21VEKVvnZ76/yBjSBN9vTUy
TcFIGfQ/CuYP+/ilyqz56+JuPhUL98wraZAnHo/2JlN7mgLXk38vAwLQz5A/erD5
qYWYg5vgloUxHiteSZfvQyWVna/YdcENEDYTxlhbJWdMcXUJfpvHQTkBCQ3Pvwfa
nu2k9fN9PmPoD6qhmTWvDCpvtqURohzeZkGsdpUH7hM33s++2t4Sb+0OMwge3m4P
GweEPnbbhN7phCCwam1XIvRjp8h9OsYx8lvKO++dxwigjvObKqnmNHQKrsyOqLCp
u6ctBPzvwuC3i20OIdLw0AI/e++0b8UGiJVlOAxsQVVglF3GfKq7DbYg7zELF8Uv
zDYysFXc3mrLp3AFD8X3BMIIxUG/8fJ6x5mdzDM9p9w9h/yO3+2yiPS5iBUCKrWu
XjDs/KerLMCe3QgJvw2cVt39Q2yi0cnjO5vngHBQvwT3g9X34IRNFGzmVzkqcZOz
9+rQyIahnHZg5KJSTlzFDzq9lUmsSqlydNHm8pTcPlgVJFBktFw08uOBBEcRxOYL
quhqT1T9iVHbc13LW4fV5EXkWwE3w/BPRk68prTJaRuDjfeicM38I0qIOeR9bpJ7
q/43LOizkCWLXtzszh7RZrPoCceUHfHBkIg19kHrfFZBTbuRpS8CEkvU+Dy38geq
/eTnuFZZ1ftgEDawV/+D4LSkx+di3zJbu1j4U6hH6VhxnYGAZhhwN3xxeFsVducR
gbEQPWtnrFqk7Ygp9246+dffLl7QZ4sHObJDIHzUmpMWclTgYjY7idRXmCxPhk9T
9gLeNT+VlN43Ux7K7nPMwLBIsb9sisuqDjEu/Gz8ogg2f/szuUzFtbMYkdhO+3Sy
swp2T5jDCVh1M29BfvAESbimU16nhofKQX2mB9Z3wsWr+6oOoGN2NeGNtrJHBoVa
N4zuIBijrTaVekkQmkgebt3afZoAYCeM9bGMtsrfd14q7Pw0hCDJn0Wo5vz+XKEw
WSIBQjaZTKQKhfLRa42T+rhGjtpcMN5rS50UoyVveKTyuVmbto+B+/iMVKiBshjO
+JwWqfAwQviPCXFQhqZw9rwSNB9BmRn4Jwj9hREWHHDoATg/TxgIbPs4qVMFxy/2
ZkHXh5z2UhQmK4zl7/kRc5EmXvAzsr75f6VQz4T4C3zbSbu4n0xQAdalorWRMa86
dKMzHn++7xIZZLLk7501F0ixlZKQIPIqvyDm2wtEtd5iUkDpYRN27OSEm/XBLmUK
okD6q5Q7JMMKZUpjVDTHi7pnISFzOcWnslg2oFA/FMyC7wvVyVOWMYHcG2tOSeSV
IBdM2vpjUTKwIArGSjB14w3j2w/0iS6t34h9XO2nVogsfoPz0iSs5CJBjszJhWR/
fxDkWsDXp+yLOLbopd2WaeETRAbLM547ME43Oh0RZSHGj8Udb0MK+s1Kr4t654Vf
vxudrMdyMx3rEqrq0W0FgfBX+nQCqlfIIA/deTnwBQqImMeUHsF6cUNBM6O6W+s4
tHMyBrm/NffDMRsc8ZBOjL3GAakcoi4YqLIhDLSKncMMk2dZTBZhtEjA18NYeofi
whm/svJCRI3vJ210M1vILdCfH440xzs0QNjiYDENQiFl8XLnVRn/WvrZQ1u3SAx5
OhnqL46IEcZAcaSBpZvLpJmVXzpg2BjCJk4/Zi5k0dWEYVwHqfmtlX6ei80DYrEX
XFCT6FSQuNLgXbTK6p5Yw6v49UTYMswT1RDOEnzppTGmnYPIZs8gKQ3shAPrS1OO
5OVAgc6ePWEfgqIdbYpQSy/TRln2ybFx4Cq/rgieeFWCwaqiEr24KcaoolesJ6FX
DxgzCBZ405FdwAVlgtKH0me/1B3k4aZ6k+6jPYwQLHcdxZ2bvBF/xvh7UF09dely
S8LePfbQns5frHyvSnJcuPtLsNJQ5Xyk3Nqm04aIlEyYKBJLQKARpjBxBgKTjOZO
3e3dIyUFR4mfvA8R0oSJ9rAet4i93GMQsEDaKk8Ta+MQLUXIFKDW3uinUT3JSjbB
tw9VID0WHLAfhnFzyA2ehsonrqOZsdtr/NPYxmjGSnyU36L3GSf2QovrJ7920zqv
hKi/5BSX7dzRR3Ba69JELlKMBnq9xgT7IRSxWJyRqNrQB1i5+8qr3/oV55f2UKhC
NBSdFbaHU8T32FY5AuaRV4jV++Ns899SugqDyL/4RTpTBbRNADCITs5u/vzPVe3v
v1+35bpQ74Qh8wS/m5UZAZ8lvBIGeMRMQ4hefZxJxIX5ECdh0d6MLZwjuEQhxSex
VYtyP7dEGjzoggGRjyvmJuPEMlZNaii+6VhoM/tlG3h+xFiix0o7sKwgPTIvDqgd
FeWTwDH7nQ2rdU+6AjWi40mBTFqAELT8R4tsO+KRUElZqZBGuLocC4V8EZnjTK7k
GkVmbyMnNOuqP8NMHZt/ia7jYuy9dK55KpVev8r1GW9RJZG1BdMbmEqgCSUHDRtk
IBmsDm9ZLHKki8dKGbvca2tSu0cFEQ+zv8ZUgrwb/7j7SFggByAsSUgV+S866+nq
PtWk3JyalEfbEhK02XPb1sevWOzLk9VmjU8EKkUk2jdi/9lpFZ6iTkl27edliCVP
f9q/QYeNz+eaWezDaLFOcxGCk0+EL2cLhJsYQ7Vu2j2b0idl36H4cttBMmEerZmJ
Qf0Iyiot/BUFfVjfi2SDwI9nAeb+hV3Cu+qMFTdF3SWGQhnAa5xlpsGtpUowil6k
CpOX5Hmle6lZrnI9NQwUPfKkyPPf4emU8/ipkSN71Xu551miMcaAWlwcFwbVORni
ULec5mg5hUH7o2abMqEfKBhPnRAqaWkDe2Vxv0Ja9sPV5fGew15UoyKZgNS0CBci
aQ71m0Xgy1ARwMY188OiTnQdU7o0Mc/nwfRr0ei0k7RBjjtsopMSEXwHV0zErPoi
DjfQwxu7MwgT1w4IwsTa6y8VppP+gpG9uwMw6sSMcFMh8VfBkNgaSMovQ40CwCsX
dU4IeKa4vQsDqc8hDaoRYOfq5S6/SHjL1E8vCi/O+GXdSlGWpSzgrLxabJh7p4/p
Z2CDNOIgq0YqbxYiGMUegQC9fKWWKxUqII7bb1sDFO7sKikEGEAoiyoP5s8kILF3
T7fuSEP+UOgZtN2220bYS6tCBt4P4Gtvovm+exTSg4PrxeoKLjE/87RLwQ3tT8vA
v3sHadCePxatG2tb+W9h+9XFQsgM0UpHPFfRrCHNszABrpwQTjcL1TWXMXP92Dmy
+jODqgOnF+147bLv6CLpSkwqysVVjBHcWbvdT66hvwwNaeoEwxIjsvVYDHcerFBb
2NnyDdpLhsIw4LHrtt5KUvbebZz1y34yta5rhIrezvHt4Pf+V+++3Txa28C6e8GY
FhCVTFIcjX+xJtt5lzlKy1zzCjSPtU/lwNLwNVGM2w0R9OgqBBgncmnlxF/FfEON
xe8TUyXaZLONQjFMSOh2Qq68rYdG3sSs+W//jHWiW2enG5WI6nKswhaGz8VrN7Tf
yL8d/Og/Oy6IRDHZl2cxaClGnsJHXcPi0AjcqZY0g5UlR7MFNdLOCwpE5SzutINj
zj3bkUES/C4njqdIv/3VZJxQCWmsd+JR6kt51Iat9gm8jhbk43DVoFNBXRFckLxi
4eVWmAOljGfNNPTVjYX/kzO/FDKWWiO8dHN4udvjSwxSQBzq73BzEM6VWrYyYPsq
TwXQeqFkYPJOeOABYb8KMT4hVK1ZkW7qakWIAhSSSMs/97KLhiCKBZKJzYzo5M0x
jgcHNuisaGm6ohGqHjtWD3UGZ4EEax4J+bgKoLqbTseBeLGWXymR437NehoWdvnV
q/qxSlyi8WxGzvvAMvPx3c8UloW0GCf3MBhi4ePL3LKufr36rJiyNFlaWRN16rSn
PP1OrBMh3OzYRBzhyag1uUStXhivZND3iAjeIVXTTPfynHZUB0Gl/dHMVeH5FAWI
n29crqSZyq8wPYspFV463zl/586J3ZGivnUU9j93bjA5mzGsNGIRM+IM92/UKKLF
a2UKeUwH1TxLmVh2peV6YxZfq05wxNjSjMdNIJkT2kFurSogCc6t6qbC5dsGaZ+G
DiYstjfUj+iHlWxTS7j9MMBpzL2+MkIcHAN1swuXV09cSpr+j8QdUspOj+/1g7TL
Vcf8lrVhnHCL3wSE7pjat9eMtHyD+JCPU7q0QObYoxf20ESGAwtpCkVNTa3kxVWN
498/400uSMw9JSl7L+8E2QS6+fT817KZn4c/+zIIaJPTTD77dG4LUXtGOadlJaYC
hXOLykg3nhMMqeru+nhXR/wVxm56XpDRd+DFNvnfnVdMGX0DayueHUSGuun37/JS
jnc3tZL4CK6p8OJBDlWWiONoGRbhDSwbf2J9l3zaq4ozynu4bjCOcnwJJfx7lQBU
2GyeVh5orGg5PXyS+B1h8hMo9YH3JA1eD9VBaD95rejy4366ULjUWTR3zzfpgxaC
sKgwlGpkfCsyG/eLeK/ov8uNf9OPq1i7WxtqfWS2d0tawKYm6Bv/KA7uGpMpxTmb
/lKeyf2orAaCiLIF3I+DLf0ijQWDa3ukDRn8EYGWvTWKVyOmwLQfph721vmfBMxy
QqSITrrVvFNTA/Wk9N9ykq92NHw9nCCtXi1KmVC3d33//mEZhwLwQTrAjOfDEdBT
Mworo2AZpB/9aBr2NfGLMVlF17syQAPSABRe+SGl8bcjgdFeaLKywESxoVSMZSas
gkcs64FylswI297jK4WClS8rNCIZFP2P7rFRgSc5iNo0JagZAgUksDZHQeoIFvNz
LLyl8OP3D/7ucgWQm6O6RzMEIdR1ZnmEZLpE1PT4/D+E1wNDutbjeRXydiRslXw3
QRRfWyJ3ImkEXgUcgroNL9E6lbk83yP/mvuhTFrmCAUc1AID3cAhh829Q005dFDq
g2r66wegoyFtrHACTFDr6f19OMXQQf+5gt6BHvb/xURigOoTxZH6F8RJKVySy7eJ
1erPsyrbXjLUutbBmUCHrRJrTVCnZuvF/f3cXPENQNhPMkmMJpwJO2prrp5GX/eg
u5J7WvqYjC3sAJWhEuaazBrmXXfFjALOQ0LBkch5jnnNzJhVufFEKZBiWf3RmaFv
oFs3M2P5BAHGNUQT2oe++C6Nlf6cYDZSxYfZzuDpRJ6yQwMOxYgn/Bvt7gNTo79U
FmLolPDwVE8SkP+QijMCpD2Ld++hL8r4OVcbZGMq6iAD/EtQTuJ4tKXc4BAlHraM
QFc8d27Ab55Tfl15LnPOJjTF9Cxc4d7819oJOM84E+qUuKtSr5gIuwHaPGxp5NaN
qOvF7RVz1WEenMZdz4Z4QrtzT+EZQ96XaGvYaC5LYTodTBCKYFXlUupBUkzG8CQu
nz+1JNgv+Je3uWD8ldudsYQ9NJldD1XHsknaSo6TlHrHBedrfMfz+ksbLacpu6nl
D01x0ZOnHatUlUGnAktWs947GbnN9eVA+/wELWcozogpX/KhPnuOei9YaTvQYNvW
CdIYZyD4GtrLkAw4TLMXCrNAUFP2w/vorXvWoabFF6CJuPfW6p+JEM0RQ4Qq7XYN
7dDUqqinIWFqqgVj8ODBWrmKacxYjdvN/1tMkADRTHV+lAh/tTOoMmDqmoNb0Ane
p5ZWVwMvxlxRu+Pe31E3LX+Ug/NEfMu6kbb1SduEOb8vBOa0E+D5cRiG09iB0E8H
mxQJSHDH+pYP9jt3i8phNQO2Y0zIj+gzCAehGqtMspmRp3mMHdYBgOlS4AN0EBa/
t1YPDnZ95PDaNZ6L5ct88QGJbHffp1XnTVO1fSVp8xl6SSn7Jdpi/4U5+RYdoj/Q
Rj/1K9Q494iLXudUvEKNIq2skjLxASD14cDmycDQD5NjEQKR282jMZudY4jElUKJ
Vgwn0m4mDdJTTIpXytqcMRZ6b9cWIavsDW3PoRdglo5lzcCYnVQJR1dmuUExoqka
6fNIXS0NVtQyCd+9h22q1coFfJQmU1hupytiranxaWZJIkYc7nHFCRCR92c9QZY4
Y6YmRTVA8Rjqg5oRVRWKgTuZYT4kJNHFUx4+yookUrgZGGNvp3HNW/b08SbG3Wrr
uXuFuMAdwk5DU4zKs8owhtFAZI0uUm/XMfv0FbDC/zFzpJuHhHXlszBx8n37RGUs
N0yUyN7dEonpRWuvxRi64AvQ3I8M+GT9tNBKP4EMlfLd7TM+69GIgkmuodsTmbAb
7PPmDNIRJU0K/K2OeT5Q10LM7Rvad4AHZfKJzjm5H9OC7nh2MuiQ3VEipLJp9l+n
XdtvZLqyMzGY2zzwrcWZjfOCpTVNHuug3gwBed5rgGft1SPy1+umOEEorX/achny
lkZqYXoHIzU6Ucc3tBBw6HAv6m4kjktohNZQwgbPHuu7Md1LCPz61m8/7kJ1K3sE
ITTBEW0SRaG7voeHPvQwr4C4XoYPJ/+GgDP0Z0ry+kMM9N12l6SJGNOSvKLxzfnX
2XHV0ED3GU19GOPqi6uSI7jlsb7+d/ZDd018mfQxOQ6wMUXFBn2bSgAxt24trQja
gW8p5dshD5QUXOy36o9sv7LyQVr5mj5Z7+VweCiO8fBkHPDbwyyyR2cjOmBD+/jg
awYRFcWWoNP/UXHYLSZub9KaYOJlVGPl9hqzpJPWCItgLqX+Dtwwd5LG03o7wUWN
i7b4nwUE2rQSHDMKb1uj7sB+LFInddIQHt9+feivTeWq3guc771h2D2/9rFAhlAk
9IU73MBtl0L19BeJyu74967pFugA70Fx5sbel6eA0Zn9G1eINl+ab6Xs/Xaa3KI+
AsrFXwVFz6yrf62zXs3zY1SlApz4Iwj5yrwOXMG0eONGkysNMNab4hzFDjJB6Dqz
GXqb/7a7wPRntqkq3HbK76z6aXNiOLoPRbEUgKP2ezJNko/h4Tk04oSdciSF+o7I
TBwJomEMAd3c6RFMNKIvhzzdXHevdNJ98vi6qLSRiXsxvOxfHjgKrQfkiTkKnU9c
d9ZX18w4SujgxdP2mRrxG3W1c3Hx6LDJbMRaWoAUiyxIK9mdP6KU2Ivn5zx2s9Ef
+gvJE637st7G2mCDm1TEi1z3o1VdBGzb2x5XsF0+flVSjZSTgcLOfH2QuENW3V0d
r0B+jF7+RffX+VhNtv9kQlFEi3gcZet0QN/nRVNevye2sXKchcRrUx76E/TxWj6k
mqVVrhWrMfHCV3wuBEYf2opYSfDOoL4nN3EPEG67DJ7uYOH16Dqd32GbJWT3kHXw
RGxdOsjO8nQmsUlOFg0BUXMjZE+eMX76Jhyzym7Scz+TSk9IusbD/PTQk8ySdX7g
ZeoahiCFf1s+tTxfIt/BNk4WV16Zx5PkL5MrL8SI/uwWYs6DxUf8rkvXZ3D10Gv7
vO5ab6LldAL5godN+GRJwQChz4TanmlklnqBdeVM3SRKYx5LJ+Ya+C1mHPW0ysCH
GUU+/3p+DwAVS+eENtePICHcRrUNPQQDq1vHP6TT7+I+Fz4foEMHTLvc5AMoQ68m
VNf09Sehl5IJqAPoBaLcXbyZsfIx69OoWbZsMf9vTiglErVcovAN3kIuzjm8DCMn
5QJq/qPnj4xtqdKgbLjxgyrYIhha2rapYYDuWPyRHnRvG/mAxKG7TMSV6yE32fSg
Q+ryEa7uMEYTEfMu3KYTRBb7affoyQeH4kRKBVBgjbe22Kf1v8gOl/OFLej/Efrt
OqbGDRri9llOcZVoHcX7ZKVusmSeiZAyK7eHM2qso+3Ye/Aj4iR6zxILDl9ZCFPo
uhd9c4ds9fwnNFDVgh8W7/nS3FpndlWdkMzBTGE1mBLDEhx7ZrCBDbR+1/k+ox4O
qxt7RhflBwEtNGwe3Ppm28YfNjVgy9jt5IQI0x8KyHQQbAZWDbAr+nZnDjjwEd6W
fSM7OjYwM69nnO8TXlQDCcFR+LkaBGFjHi/P8RiIFy+rqHJlmh6OQHEeTJXO3fUV
OuuccQIP00G2JwgaoqecrrHrQSAFaOEbes1Mr87WUdDTmz0eegJ3TLZzvztrp++G
qqrtVTnRFh95zmJojvPcz6jgli+C54DIXTXBiIq+n54PWs1IrpGYY2Hi8ciTTUyI
O3C668KcF3E32Ag8T7DlRa9BtunA9y7CTRXr/1IYaQkuqDRKrCCVnZoa4l7/9eZP
cGBd/2imv2/WV64kAAna1KUDm11PEwCfGbyci1YrRJe6Qibyei1GcQ1kjPbA0rWm
VjDOwUj97IaO8wBvyC8SCognc0t8ky0qDSKt5I4OEWe0sOGNFFWlJFr5BTj1WVAp
O7807UW857TwGKit9WbvVSYeYlgAMXnX2VMYg64A3GTPwDtV2MO73+VuHbouwzj/
Nbvf9+Lr541ituAiAy2X+7BF+M6C7KmstsjM3bCbGnJzkZRHH5SYAcWha4dW0ZRH
K8r526oWlN/lsjk+lwcpxjDAddib+UiZgp+FtLuhzEbY0UaUeK6sMP/Z4f5hw1un
3pWO7DsdNllZf8Lb1OvqABs+4GR41/+6P0iLX/neTKv8AwR/0Z19GsCjW4sCFrtP
tdEJEZUoxHbS4l5lCDQGi5JrhZNpegSpM9oTMr1KuXzoXmNHKWVbwpJGtDLHTER7
7O8R6yLF/fEIc0+nC+0u1WGIm598pyPx8rIDn4GEjbvcOMNw29UhPD3v184tDeKv
Gs+rfyc+9CHe3C6t7XSVFpyMErNLZx8MkfXtCYDu/qu+4SRB4usXCA/iMuLs8s/H
2454fjnMjc61e2UxAEBQE1v9+JEsAkA+XvQPQvHJFY75pFyiu29yxMZaMG+fbkwy
UZqrKk0dUGr7o0qpPaVReCCCWglJgGMBKPmWpXBXNC6YcWlmbJPERX/NIFR9XtkY
EkRUJM9z/88p8Izx3RLOHy+8b7iV9UKD/f1Qkh1dIBzd3pH2N6i8HaGpg67PXkOS
2kHI+gW0qHg+vq1ex5+h8JRqk13JcjhApvu2odpNtrI0iDxfn4l8H5VCGph9cSKY
+0LUH2EPDJcUbkrBek5MXPcVIFCiLheP6U30Mpyxqq6Pok4hDKDMz6SjFNEwRk85
JzXtKR8uCJp2zz42QBRdBX7LU3hN48RlSzZUjdYomvAMGthYd3XjDidKOzISYYZs
0RnRZrbX8kzmqQvBeEdM3D0Lac9uGhy5TKTEeULH90o4z1UCl/SNujmxtfW9F9Kq
REE5O/PUhaC9g831RG+J0H7ghNpSRHdSM5CyV+X4fp21U74PfIO4eXffioVmP7U/
1nsxU64lMg2adxH9eRqfYTPVt+vqT/9bNIjqIcztzx8Y3CvC0d0L3ldkHPCwV1z1
bDtBT6Ycs7Jufeo6td5i6IaMKOd8OfSDj3K+pubFoyM0KRP0tJ4mQjQ2daTDH3px
75y+37+LI7O/sysYV6qHVQUbkJizQiplQlhRVT/YbFusr//jxN8R7cloJEzn3QWd
7z9QElKmP93SfkDInidyCvmAYMXy3wyIPfppSIzuJrnrgcDSKBCagSa8VVlRmZM2
TN3cuKaly2FB98KqOzU2bg6HNJuELEwlfCLou7AATVyegTvx01Ie1l8Taseydhey
guie2m8vTVl7oIWgw/FtvdQqxrUqvBiz3OS7QKuXRpy6bpOhw+KGvFN08vGz6RsI
AAZ8bfs0Tji4ZS/KmpDkGHJFsSxf688kEwQIVgJzU1Wxq/myqcDF34otig1JZr9r
uty0ngP1j7ArNzpAyBdvQiKb/PyRiHjBTHz504r/vmrv4TOcfc9piDiquyiEumNn
sxHajfXjteJIc1aw9/rdzAJV3r5cIHBRNRKnDok7gCxIc9VLIWPvjqL3DKkzOWXf
5KnWyO4ZOkZ0B8GBa5EVbVILHKdleewcP/nMRifT0UZ3z/Z5e6LiFbdAUqYSdDsx
TPJCqCIzF/lMV83y8g+sQ942Rg3QBBvXGPoM7hBkQxW1IyiBk9Ls092yeFXcqTNx
9Y0fZ+fHPnzxOGpjTf7czHfnflt/RUrKPa9VK4OL0MLj+ax9YIf7pJ+ql84dVjsq
/Dd8BrXWZ1MUXMTyRiyg6BONlxD6QnQgJz11g2uJLU/roQ4a6ApZaMWFJrTNNm1X
MdWpDpjs/ZWtArmIUFSdWqWLsE1oRDs4iG3GtuiPtMzwPcXVRFJwB43rQcXKC5ut
1vXaCwUVUQLJdEFy9B/3HHoqNSkzJb4tdFsCzDuDoLA0fKmn+x16OKGX5BwKGxQ8
AVCFBs0PPag8iyAMukmK6kBp4tTaKiRD5V5K8vQaxEN4XI+VrFjFNRaHUam2LF6e
6G1anI5ZfCyM+w8jBSPyllzUCngNvTw5kbcmEXXfj/t81iVU7bbTfx94EmF1W74G
MkmX3urf78+AhxYvVt1VpEkdt9Io7iuQiOs2zaIxHsBs/YI/jwG6/XxO1RlCClqk
hiBSs6/i9bQB2+DWE3d1TW0uu6eBRzc0RCWuKGlJvlIhwcJr3tqQqkUZ9F5z3FiE
yg25Ou81B+m8haggZtATxuPY71ed4XfbGhODn9fOyVG/KtRNgiLoA1Vj9etzR+b5
HmIfGwZXUOs1NDd6WRMNnumxqrq1NVO3pUkB26jE5M4DUk2GVWpM5qpPEG7JKRe9
64YRlAfcOa+Z1Pvfuwbn9nASkWvSXdFzNhMUY/hfsfPZ0TUFKmDzYUrCJS3Wpjr8
PNnF62O2nxxMNMroLU+3BIkqRmyxS+AGlyHprB2F76pYORJ7l09XJlJRq9UgNkMW
iekvJSf7KUhglebgp4cNB0wdhn+4O6iSUnan196lfq4aqElVQ0SXa4Xbhh+Gou77
dvBhVvOTJeQagbfd++Fh2p2d0u5ORZRhH0eOkoZHKb68o2PESWo6LuYJi3RGNTij
kXuM4RDy8EFrmOSWS2u7ZEW9ENgcDhDCiA3Gzm+c7oHqiluZs9O+wl6BWTagXbu+
4+FezHHK8WaYegA7iyNvwnDRoPeReltZZEMqiFoHzenK6NXNaH64i2+1b8cqMZY8
0Q2k4ObksK/34m52rdQgTpdgcmP0VCr8bKLT5mX1O+BtmtDDl2Yu72PLweKL6HZE
Po81D0EF8dGDtmGbmdewsFq3tc124A1Rhf81ztMmfCDu0nLoYAwMTugg0ivldLi1
RV8W3xL+gUmB2pv/8xCNH5VzHvyfn+OGg1M10Ew82+aWDZWng2oDf/Ek5GRRT5I/
F4bglBQaSlNgb/gWPQHuCIz30B2zJ1SX5s5d+nmzIKZ0ah059IZl1fu8AmTMbpUJ
zuhNGbSidpv7O5d3n9DhWhDeyoPouTPwBmRsp4W+RIEZHaCRbLHHmWz/0uTCa7UQ
LcJa5ywipr6WCUppyPDIwQaD5N3hXdoqwyxHS6dyGHeZ+LM9tjPglVkphJB/Z0/1
mS5rsr6FjqaLhhSGHjv0tsLaAvIk9zjiCpm2t/HjtLsOdxqNMxpJpVkxnB55IAQm
GdEe/unTH0szpNsDwMPtqTW8oHuniBAF/a7cKrM1c+WDD6aZRy0OS10BkstFkTlP
Wlh3VJap2XEEjM3JLYJoE0yIX7QVbTEqqKpeiheIV5wrbmaYT5eVzNJFSQ27px4z
2VmZFx4tb+XSwBTBmOxHT66U6pkiapta8WRK7vM4j3kbMDVrKBNngYqDe5tXVTVN
F1S2koyulMeBKOOAJNetHbjTMc63Gd/dN4FiiE//hlrMvto+mDI8C796o8MJVJoY
jfrtKf7wJJrPzWAAvJVsVFArrxD40b68FY/ZUmeeozhopFO7hSbJrvPlcxIRsqTs
RgPz9Jy+3YiYkG0//P2oISqkq9wcK79tQDSW2dY2jnqVqH+JogPTGfytVQ2zft4e
UsZz5QIgvmlsQE/6d3IgrFMTadxZQmebDcrO74I6blkWs+WvxfzPvgf2JwNbeokH
WP59W0wyXP5by8zZpyOeDJLVJc872f+yWZUAL1HZsSV1w/pY6HS2qAhxSogf2JDD
df/UNyMY7uFnJp9cgJe1aUcXdpB1yJTtclWF328x+gbRCy5sDlEEi9P5nX8wGN3c
dRXQtuCEH07V5ZtR8mEOaqbWpwWAXdqbHYBF5kVm/A0IH5zUmc0uJvGKC0lR4Ttk
YjEt0pZamgTUh2zHGRN/u5hNmwUlTNYEyeYjnOnSEWQ61mOG4paPBO47fB+BAmyx
t7TjaGYNNj2FgC7B8zHRW/tQ8alckgdtoPsl5sbt/r47pLSNcTc5TVBTVDSvS9Mx
LAHGeWVZ87FGxF/KNxWZjLuy/o+AUnPOA1DQjbva8hCH8tKX3BlPkCanXvVlResW
6qz4byd3KdoYZP/agR2iOafLqnf7RYJMFLAJDc291ZV5+crxCj6hUiuNE6Lbx6Ou
SCibaHgbKXUwuk0jFblHLcA1cy7VKrtYfhQnsz4FYZy+ue0xZSmh3YwkMWMxrLK5
8tVw1PT9p/rnrq0LCccV65nPkV3WmEielY59Z/+N1i20kB3wx+8808YjxtWaM71L
ecT/sMO1uO45igSzvMj67OIgUAFivl+oDNbinMZf1IitQhPpmpkANfpSlWxfyNE8
WZTFpExJhv44Hjm+5qh9MOwRpfS5yKrR3W9awM6O57hSQlJvJgBT6aB43tr8IWuZ
gkSwDBa02Vtedk0c2EawxTivYfhfgSxYT9IssoogLr5K9a0qZhQhPu1Bzvv00z9G
Ezsp/wExTdDOxrc1P6fi8FPPSCrUTrgDfJV8MpF6vuW1kyV2veP8/6dCsYnkND6q
26s5OGMRotRNDiuJ7MGKy3kefzpLvt9OhXnikRqSWXa715qzFwYuzBonEuGu62D1
MLY23dUPEWvdvZUpa9bhyHa7Op4RBIVbav4eySWsKRL7dIQ0/5hVugNAzuCQ9tXf
gq0F2l2hB2YipQ45LPzoLlvJ2EPBVL0zrejg7q7dJdFevJuCnxQdkL5rBvV2eWel
pl8IbdUuRC5jjBNgpgLg17kscL6LFTvglvKKKqNxEmOb8vxNp9Pe2KS6eO8rDpHH
YerRUH6yqI0VuOr6o10PNEjJevTmN8rwH4kR/loN5K8hxDBs+4N3uYMT5HsJFn8c
r8JLRcJn4jeAV6ZdgolYuAq634yI8zU+Q7jYqJPHmHHMJM93yOg7+0Qk2eKNHBSL
7OjWCLZuLl0JwY6O1R0ye5Rn8t8G+6Xj24D/jGOOJ7U2Rqw15Fp4vW26qENOPwV7
na2L6f5z9J5876zdwdPn6MBvkbOTTpG2DhW6pV1D0nflxXys5oJlqLtPNlxZ55Ex
NNzRNSLCEAYsdVyv+nNEMbQopM18Lv+xFmKES+31kZsCuZVyxeWR49OfTP1eBobC
6AgMB+VyuqoyrNTepso5PYmbOTMytQyup/KJlMikPScxxLPye/U1wgRHeMDIxomK
skvQ5P5YNJ8WKVPPqJO0HWct60hZuzskF2qyQsU1GTFTIzLlmoHRAUe7HwpdmH+C
kJ2BL4dyN2piUI+SBbHH04oLvppS4rUCofiiKCKEvzsyMY7sKEOByAG3sEj/77Gr
YYvPe7A+KkRFNxtpgWtzvhwoJIXdXm9tsjysho55g0CjtQ6n0gihfZ/DaDRetMzM
BXmXhp3seTq3DXqVixYmIeYuHIraDNdzJmEbSJljN6RixwjtBWW488IcAxB5W8lp
6szDnDzKhvFjREc2SQIfPCeJRQlsYN6Z6kCcMpIDHXtWoQc8zQE5pb9K0bH+NNJ6
NXqK+tkohx+zkYPeX/GOH6z4Ijixk0OCttSDZtCuEme3J9LGZqpL/umqQijKycBp
FTkq5WpFEpTD4fybnZZOG5VBlgMi+t3Qb2cXH7ucHXFGbFQbcmEPbZdRNuG/yEFc
6MJv2itz1OEuVo4TuXGeR/JcSHfSIJ93f/wkw1TRnY/aW0hF858qcKB0SCSLbfvZ
8XaYClIK/STEiBhAtumSE10e7ae5TBzGqhNcL63DW0AZU3IpfegeF3dgEtGKSJE4
efjtk2gZRNO+pY83NCbivzK1lL9eeuWP2FH14cMPBkvzbyR5ya2+91L4tHVmkCnq
m47Q0ifzGyxf4AU9S2DzSTxXFjweUQxKSq4+RNYkxh0joqTD7FHh0QlXPsduonWy
IN18RiVBETxggYIIN8imL8TPS3l48MWaf9BymG3eLdt8FSBg+U22rWYl4JMcelVZ
EaisTcCl9fsCdSVlERfITAq7/4wX/5Pfcoe3BnaygTg3Ka1MUV49NBR9+TodcXyK
iXJdmPjjQWQMU3v5KnK97iQ5BaG4Cskf7M0ZlFoYJf9Y/txHcKC2QwbggMpLn4IG
8TT5dq80LVeOZ5suslCEY1jxM+S+cGm35nzlmGfvXdZrAfU5GSkX6QUeEjsuPzvl
G/+U9+PNee89TAjzAH0VV3vWsP4jtY6r1aStdV4INw+mGnpENw8T3l3QHcHc0GOO
n7N9QINglz+ZdNr8tJvq3Bn0tUmBAzb2c0nJJzA+rkuqZiQfQrLT2X5nUtD1ysmj
VjuL7pp8RPCfuZL68F3/62qqCNEbfqT23p3i17nzxJdf+/4A6fkvXCQUk8xp30Ua
+sRup0Wu9xTIM8m7a5qFQwROPDdR0PGcrfDtsjvbz6ySNOeYcLvtSZ+YXteNqmrk
diIIFxxP4bwY077jENfZQwGiNn1dn0VKLe634og1/7fdqmuhnhQUnNZ62XD5q2cC
2PY+o4QpBF5jcI3VPsDhhoD1kAnyt6ppgKxs+PYc7YSWxqTsSL5PRhNEjoFQlz6l
MmrEJa6gNFNSxjNMsFG4DQKmdaZXT+fvDdDOlycMbNZ94X7Kt6srMBjNqs3GkfqU
Nt2+dzhlZGQrg51r0iwWOYLWBs7I1JuAAXC97yZU0x064umq8EzX5abjT14jhden
ZlLe7Uegz4xEjaDoTsxlo1Z4NvZWxcS3+KQDp5p3jNkqGH6NiWf8RFxw5CA3m/j/
oCvWnAaWuBVM1vyqy0u0undNQADJ/khtq3p099X1m+LfkRNsEUMAqFr7hKXukpBx
jmLl0lx4ykN33rp+msAoPfSuec7pLgZCGz+kmVPcBBu77sQXey/oUIiPxgVl87Nq
tgTjNdYoyClpCf3Zq+CEd44XbLoaZzQdOkSeau9Ci9ihnTZPJCi8VHsHaJWMn7Up
2crMxryemYahPaxInxPMYlHFj3A8qwOdR/HuvfpZufi6/pCYZiY9egL6Ruznapie
yW+3oCyz9hOYU0sFQvFCzfQLCSFjHe/vMu7ceimA1C5amMXxaz0eqPyctf68lhzc
8zFxbVDKCNTPYZOxtKZP1cH/8pGuBVP5ja82djqx5aSunDsPMvSlpSrzCDMYhXL7
FkWtbpuQMY+IHyamHh0oj3bhDXWwTPSZs3gsBbrVfUAJuWJCJrh0nFGHMR3ZZYVn
QYTR9p3lQAEohINqfmnWQvvXe9xnv6PlKPCYBlPsWQuiFQrso98M7sEuvmnvvUnH
ibzE1rU7XNp1lkleG2dKathQ59lK6xaXRTSS6Foke0Oy6e7TkUKa7XlZqC/CYdm5
vEgT+hYXM8xGjJJBzviz0fubVx2t//7EtXIk1Wo7GDlAQM4Innt6Zz3XwRBMYybs
oY4j9ZNo7ogL9zT2opPTnd+HHKtPPGUxJvrqf169BjV89b20gojXWWOYQlZ/pat0
r5Fl/DHAD8GeaRkarax8/B5bZYfyVj8AoWqEM3oarNGRoZfTavAUdEfvGfHekiu2
bQ7LpJS+LPDE9XgY9O7dae9cMPKej0G93w8vAQd9FgzlaKUovhGfq7xPMDjaqTJq
6+f0MkFa/9KRbz9EV5DKslMHeV9QWsNj2EVnvamNjD5JOQpaMWVIYxiA6ySeLt0n
9HiPqaz21LM+c++XBD2mgAwax3oI+e5FrsWV3N4NuxbI/Kp6KhQ5HplKTh7IiPsf
UiYAPge7tnP66YVypvYglD+TSukXghnSqEfX4C0i7+LF6z1F13ps3kBnR/JJELEM
PnkYET6YWR0UG2Xf4qhsWxWotDf48ws5x/HJmAxtZPRW3voWFdIutD/GdFkltvYg
Vw9h3cKBO/EuJVVp2H9+k6ljU/w26JvCXZlaIR99GJHVnUIm70kTTZYfGYEDms9T
FVJbp64l8sDprpon8HId5UQox+ImcyDCL+5zouT8FGx+RtnBGbIFZvTuX9of8uHS
OwiMj3crKm/5Z7izhGKDmHfuEwMnHn377xz70CXVhLvmsdTmjLSI9FE9nI57daqT
l1mN3m6QVWdb2iEOPAx8/SomY1GvM3jha/zGeUlXjGh4p+T5OVLAVSDrLESwjb+V
VEAiFtC8yXNuE3Q2hq2wFgPr/qJyN88WR3P6OGwTA0cnL7CEyAy5AqYRGKMGuu2v
VlpDqcLWPD0sfsW6bks7CbmYKgFxIdjH5JQeFtmEakgfROnJYAPKtwDc9+eAk1VS
WOjN9XUu6p+zjZI7L8hV5UPcFoTx0+INgPM+DnlCCO4cUxPUICUqCUmChK9WrsPW
HTcX6+gxgmbrYQDN8bahfJud1aKYtoMIXXmI/zhP15Y1fsDULNcnaAfTL9WtYQgP
q4CVOcBXZBgN4LPD7LuVs9B3DTNsuZ2L3MKHxKPJl/01K4qS38dH58B9cbPr8dn5
m0owBrgzOo2eTLPzNKBBbWwvWAAU1qYriO9oFGgHln1GMECZk6nQSvpNK5k6Gmf0
/iU6dKJZ+uDZimHI6y2hAixNCIW8WXRMHCzN6Rc6LvZRGADbXTMIqCf93G7trOGz
bfpOWdx3TuPBr2crvRuxEfzzPLNUJxvOmNWA7JWVl2Jy3EFP9ZLamSlJuImLl/nH
Z3l9+dEdZJEOD732rN5g980SDM047xa06ozBArEL+CSJ9ogoRNkNpTf6E/QxmsFJ
bXKMvydu6BQ2Cj7SDfm2OQjGiqCXzU3RxPmyqGxWUCHig1GQLIa+y6XhF6QPKimg
deQXOo7/mCkNUvHeXZMxy0VXN3JS48Fhtz7Zu5MBcSj8OKhs69c/xaM+kExT2BjJ
NUmuDI315/Qwz7FKbienWNp5NycviPfPosxnrplH9D4mphJtPzVMW8YS3bql2p15
TWSs47MbDM6MsSPnEHmg/dTo4whWd6NI5rZcq1oFBMzGuwRNp/px2RVd/cq9WTCl
bvNyDRuKVC4tTPwo+IyMQ1xHLvLt4wnET+pU1/umXyVNf02Av9n8e+sXpl7Xti8Z
6xIZ5xQ1nx7LFUOXgoYfGhRoiiUtXmf8Iwgiv6IAhXijenOK4MslMh4JdR8tWQ/o
levEQlPES1rxNQlndb09QsK5ho2TlNJjYrOesXe3uEx7W+2766nGHIv5NcbLy0Nd
+MnnemopWYGK9YOeozBroADh+lyTnLML5lEOxVFCzcdit06+Hf+Cq6CGHXar31Q/
rk102VaaNFQkoNom4NkFVcvkp9VHiW+qeIZD64k+lUoKKh8blaht+wtMb6MQlTRn
cURbCLwQTJSstpNk4juqoD6a8CgnTdtcKedPeCtsV8CK6LDisNOWqejMw0ugdS6f
Bff8ooCT2/0mfchN8hR4c1HBVOPYtAFROhpJlF4K9BVzszQlhJBcRHKWynoE6DF/
2GNsOGEbGxxQIc3qB4zraHLl4bde3581R+Z4IhPCa1GGUKdHSIuOgVRMTB3OxYZb
NUb+RmFX9gV00bXE1Tv82Z1Y6clPxW8YAOr37MhhDq9L9sCrSI+h3HC2A2C5dZUU
HJsxGYMMJ4qFO52ftbfDGFM6RPXIQxSCqnbtTE1qTUf0QsUzLcHQFAxBWuf53WWE
5X660f4fd/VeYamOfBSsZGhFn8gEyGK1BKDm+jsjSIjE3L+sTWj+npkRqTFqdDX0
MWmDrx1Pc7oLtAc+QuqGGrIDeh3/9x37dXmc0wNT4MmepefErsjMZBAVA1rh6ACG
B9aR8Wi7wn57xtxxiGRZlyNP0BKn9ZVwFWPTAqFdqhnt0QC4hPMw/JqRCd5wy837
aloSnYYgBJ18FyggIvU+d6GSRA+8F1Dz8arVyJIBo5eO5GnvrCP+0Y9bFfqEHjKz
GwtqlVZkG0B8FV16lLFEygpYF0wa6GliQLX4BuQCCIUKjKPbhKUbaC3v2k8brq+y
YPeF6MDT3s/5Lzb+jCjO6tRFNN/TlC9ULBUgQPzJXrP1LC/IyOvtiYnqsFQhn1NN
4/QjwiqVpfAeLi8cKN0UVuHKqNt88vt9IEB8u9co7UtlEXYjB5J7NKI/XqSCocpg
rLTQWC6+hfTnjscOs7AZcWOY1b0jbkE/nt5Py49NRSTIVx1NIcOC96LW8I5sUiux
FWuJ0k005pru/2RQD4f/TCxSit5a6UWgMlK/lpPELX7qbp7zxdzcqb5aTlaBD8Tt
2BSqn1TZhfrYq55vy9czq74lfVj3egq17ptaCjxDuvdt6zJHmO3utSXh5ty0hLID
t1nhnwvPqC6bfwvSidV1fDSNcuglfDTdcxOvvp9FlQeyqYn9Voeyrf1AqUf4SpGx
tjbRYz1lUnCE3q2qOipSlQNn21/qt6IQg6ipoWrp8tQMjRFBajzraQrd0OzdHm0F
bFxyIibLckT4thXjpdTEx3RfIAu+2iVB3HGSxulktD8Mta7XTk/aegpYS41e8JHV
vQw2L7UFeG3Rf4A414C8ifNukB7dXXBOZgPl47Vd3xIG8OWeAbhKeFgxH6afFIqX
JuZEMh7BGb1FfmC8tGEr47oLOMjXQmeMRk5iOhy1wIRxVF42KKTW4cmO2as5G4+4
9aIKVKIk2bME052KErBE6UMHlXFgD4IaN8wZEhDu4CEOsx9pAXJSN0sSnEwpYS0e
vsK2oN/etzDpOMEFqq6PL6pyNuJnh0xAEabELXGV82sJ4fkHUb5LbUYwvQQRKBXV
raCHRr8cy455W5EWV6yTJWiYRFvjqx12LHRkd5Os0NbznPcQANd1ybuuns3F2VWe
zKuPReCiftMqIdVb6/yDFWztRbnfqEm6/umz20zX0xclY2serygEq8mmUxFmWgh7
mwOvQVqL2miNpgClYpS0PW5V+lIb7paUwXO7wJ/LJ/FUJWEvyx45KbyFf30mk7nu
ECg0YvZHsU5Y93mEtssJF8E0A6ZUfXd1iq/d96zulr/iHLPYbS38L+yT2hFRURuQ
Zvnzg4SRxANbdc8j6vVdbl8B1uHaKOpEcsTxglnaGuBX9eqervUzmjw9/uEw0isg
OK3NmGWBxSsHP9wm1Sn/uQ+gsgEF2hFGwcl6B3I1Su6SJLsH1mCbklQ+fcsNOuWj
TFJqFK7AuuzIIIO4JhPvKbijt6GM0S9G9lKLmoJd7qRY4jD3flXxVk1HgGIsO57E
4a8YHAn/ngTAtwS5Dlms+1sqO+VNdqBtNWQ7964D+/L4sYF9vNuccwU30Yxdgxdv
WVG+CI7AQ5fhEsX5wJ8PTuwBbITQUrlPtsTRvq1MXIB5iBUOndQpukxFgX7VLMrr
fKHE80NdeRNRwrAmcdMEetBCrNmke86IGyoVj0TceWHl9pb5SGASBvr6EzC3rGXi
lmOd69NLq4eTWzb9UH/ehmJSjAouH+V2Np3NjpFVXyJcRETGmvoJ/CzZjMkIlVCK
D+P+lW7tLTwGXLm1Le1e1MnjILB4LkmaGIYS717c4dylz+NEszEpGTnioRf2VOsR
uL4wOfE51ZK2jnBMkoeGp5OzQVgVOZXP25gkfBl+1Pe8SDCgK4W1gPWHMhwMXHX9
6Wqmebig2Q6TzBvOibeOhuB0cTfxcV7tDDLk9Yagwexq1jP00t2M05tAbxnsAs1z
eW9BscgGzMCOhNQupn/iAtNeDRENQdsY537y457mPAT0sax8iQN81iu5J/zt9cql
hn96njN5hy7fw0zuMYZ2d472HQ8iI/A/pAZTUQoVPOGcyamTvpPfNk/vZu1JFl4o
4aT5H9PIhPkjKzgKwAxJk59rq9H/sT+vy9efOC2X0PRuT0Hyt729HC6c4Td04dxz
RNTfSan2dgL3ZVP8iLqP4OqlPPCKCms59hkljaHWz6DH7VaeUpy/EgPRLSIfo60u
O+kXqMYX/hoT1Qv6PjqRojI+qAfljqSEG3F/+Y1afaZaMYU5QZVF4HGxaTYWENA+
m8FE9gwTv9Z2/swvZiuU3qA7/FVYHv8U8xgA5iaoeqiJt/5N3bjz3L+r5y7xtPGB
eR8BCQY/SOs0aAqUBP19Mw7yGOSCAv75DGMor2eyYpWDAKy1c+As6Xe2/xqM6aAV
YCr6dy37BhE2GnKpEWt3oMRDP9iiIpDNlmQKeP3NNJji2ZnnKdVNM7kfO9I7xTqy
/X6RH6gbR5nArCgw4mGDG3IdJoeCgZ6Bm2e3M5EVL20bOODnmGJiXsXqhVUjq2PF
c9j9YhCg+9XVnZZEVh3nkNJqiRDilIIShGL9ABitbEMsoar96RGAHQohXXvd7AoD
fHECSTx4l2hX+m2l5BRdmKzaOixGjxH7fTY3qQ5apJ0lR6MGXHoVisOSck6GdHLD
jDvEAgb/dCeqVMGFRFXnx5DsGo6LkhmxprznI6LQQAf3lDNYW2aJ716Fm8LItWSA
ijFMpZBdinSzrxMUn4VKSDL7u+8fNktK/DthIXdhlkS2jspxtWhoZV2+SirACZS3
2Slkg+ljGGrQXwEcyp2KvTB5jPnEV5/ggbtI8pexjfbH2R4I4skPX9/WjEkKaejF
woDj8yUZgY2qrhGrLfYhqZgeSlIKFvr9xNE0ThPImwDlQNwrsdi3badX2ldlUQT5
dTwseG2ifVxCVLOir5kzyUnWrHuGrL0d5igzLZ/QJierxTIsG4lgqqbwMtgJfrqZ
IT7DcWZdS2EK6FhtJtm+N1Zbz2rqFXLq+pX8ktd/5mBYIQ2l7ZwF9XWWcJu8NrZa
xn1cgR3BDR3Tu0q0RxTYOpIeaCP0gOWovITktiozk0wYPm3tEzv1b3nBpgFItSjm
XpOxS2BDsw8a6fvgjUXGGY8QPGVYWPzAOmbQFC1PLCDOqKYS+gA4ZDqHbv34nt6J
mWcLq+23W9HItuAcRgBK0PWOyjIGupRaStfBlhrsx6ePjhXBJSW6T1q2LlDZlqw9
DqC61lmkRaTLP7A0MqU32m3Wtn9flx2eSmoYQ2YNiF3ucOXT/sreTSmi/udE9Fm0
8wVf7oIJHswKI8pb+6ApaU5aeaSb3PkRkN42gVS8lcMKtIGiF3cfy5j4rZobQAcj
5NdZyTb+Yq1XvGtMC1wmXRzYTR0QVb+E4Il7QiIskEoEVqtIvjqqZo8ICrqb/1Dk
DiirWaG06yZi2v+RpIzkrS5Sp+s3byb0sm0Ochlw/m9alVV9D/9ZNVJVlEXh6fHe
hMVv/qjUh0rpduqgZfzMuHiKeguth3kbzZcBmK28o3WVwVEIOK9ulIluWdq6l/x+
YkOvIhh1sqMJ6ghxSuASvN8eRNdwh/46L3sOENOpwyJEjc4DTddX1Rr5SGNu/abD
a0ehlHfzojf7TRiXvJPf+cQWyuaD/L3IQj67eOegprqToUCTcb/UEfevDfZX7X+h
wxlgJigQj+IaWwSryZLnXHrLAQ98SZTfKPSWrzlBqrF53FTwJC1hvyEaaqN81yxG
nKVB2RFcM1Hz/N+U+ejAXVNixKddXPeO+adEJqfFPATTfIbSsVvnF5RbYdF5XCVV
jYQtoZnsclftHwMEUnk2VWZL4Jn1N0KQXu28sxpzzplk8MPXru2t1bNE9cRdKzeK
YI6AAM7lzSQ4sOkg1YroE3a7QE99jm19AOFx+11FxJps+n/KOrmwjujSlPP8Zep7
o0GzvLzOREDfqhlsT7j0qPcJYwOuRIDdOrJJyyR/7JcMtjklh/eimGi4tYQdm4du
lZjVEUBoqqB3zPegsKXWkCP/DhGXam9DTAu+l9VZbcvqB3aCi1sY3TSidBL2xS+d
v8LrclZD/7zOdXh88QElc8XN7QN4BlBnCipLCcTCE3YQOG8tI0R3xWPjN+0hE/4M
0f11dmdnMfpT7n7COEgotZkTYyjhaIXRr+FBzwgi3WE9+2b26q16adgUWkx3P5XU
7bflIxw8u2pTccv+YmVAeJ28X5XhzWqZt8Uo1SjzGU2kMx1TszLXQcx/D9g65PzB
wlEZmCsfDBgQgbksSiSQdnI/HRhZhFJIjfwpPZez4qX0JHZ20YgLupXHtWKZc1ES
ZAlb/OvMf3bx+Kvyv2pzo3oS2+5SmD3pj9Av/6fAbVUfY9nyvHMSCW/rhwVSKqaY
2fEIcKWpAk91kY++du1ac0T0o3URr8Uig5iRJN9FHXsQ0t+p4+3tYEINjr8w1Zg2
9seTXATF/iEzDTlJLXdza2QGkHLCn8FEb3kAk+VsHFu9eIQSCbMgtSbtCPjxInj+
fA9sD6Ow4mYEFiPKBRWed81bZPU4DA9NFaccGAVQ8+gqf6fmWJHrdi5vS6o5FTNH
76WlpGsFZ3gZ/AJp8kEvmnUKMgPbpeFXzNF4JRCYh4xu9qExpSMkEiKKelDHurdI
T9zTgp2yb58fW1hq6IIzES71YKQh931IWWiJ5dY/9Tydk24YOlCDEOMCuagOc3Hk
Vyz05ZMaVYKLop7hggDGEutdw0DiVsS7Y2wjpgFPf/Jnd3+9hLdL9uft6oHC1fOB
fMMHFYA3edrlu2OwSMGIt6entDyqxiJ4u8HiiF+Ns1PAlP6Wu5LUEUqyyDtwD9ZG
+nJAh9HXoAfjNVDFiDTNyzi86RXruHPdySj8oRgWlGdakUPL4Sbv+d0cMt5mHP4u
x6WQXfA4AhX4KKzy9mvA1qLE6BTRO4qqUObbkbncTN6a8B8I6ul262VwRcuosP8N
pDtMZsFXJ70zhTeNrK7GjBlV7I/D+x1T2TOkmk17gOvhcQ4zG/5GyujkgREnt+AB
9b8Osu+GXqScVRBJSgq7TN4D0fOyEdp8cbHQHXPl6FJW6w3D2QuftPmGE9edOJce
5PDMKrdRQpEE3w2c9hWvhLGhqCU8xNPRDzkflbC/e3/YFHoaQXTUXfWAxa7tNjMA
9G77l8IuyfFFXFdutULuX4QJvH5LWWTO02vyLE88bNJ9dW+35u0yX9ERjk+GgsYK
DTjLhrRvmUwiMSuWoVNU8DrGhSku9mfBTrTkj9ONe93Fql2QcOxvivjWxV3lWU6S
jQzTgRkfnTO6WzZDvqmvWzkfpmeKkwlEIPYXORsj7rgEOZ+nTYzl2aY6wrk7SX5a
HBE82FaznJmLHbcglEg1GCWvn9sXCKs0JWibqOEA15zD5uEoxyiPRGtbI77F4RLl
lgCz/yZ1jc4Fn6QSJCpgZ+7sr2QnujjxBx8KNEajVjuZ+PZXzg9+rPFtXkO1U6d5
69LqKcLaAzqEKW7dFv6OvLsDxFqFDCPcn3ZCM58AUXinmbAN66xZ/ijOYG1syGCi
QabOQiHASjUFb6zS/2OKdVRv00K015czZ+e2GwiBLU7+e4kS0Q57egFkY6nD1mrU
iJVapY+KR3v05knTtIWlh5nNLxPI+udP/32vTvYfcojX+ZE3TQywd8yImUZl7Ndz
3SqiWGDO1lNPMa/WBE7zSakqoaXqY6Een31iTj+mwAErSuQRa8W9oHeaZffTwZfy
7UzaImOFTZm1BVqOPGNZ/gdDmu+YZi3XFG5u5QL75UUnmbtDS6/mynihH4/rWHqp
CKPIKNQp1m88t7NJF/kSMs5llVVT11lgJBKqf4LKGRIlrKGH2wdq4FkAZ5OWjcp9
ieforpb/nE3uYrVW5LP5Lcp3v5/or5/fzsTmMKTqoh/2GOabLzOQ5OkGJnU0Kyzp
RjM1z0bAAtT559JvVF0PuqlbXyT+vy32/HhCIVvsgsUnW34vYMEdE//KL7iXB0dV
NxctNvgTUywd+9EBj2oOji1J8DHt3AlfY/8iHD1ZOkE2FgMG7/lcNonA0xDzPB3F
q7TjWgYWOfzeJBweEhXoHWrAMQvLBQ/exXfMHObWl7IDxKQRdsfZGk+6woXDkpc3
x4DoTAPdiaEyhQD7aHs719cNCr6QZNx02dgC+YlxKn8O1PwMVXl4adjQs5C6FDa9
MOCUa0dTg5o1SG45YK/aRAWG6VvEGPpxPbKLhTicPT5tBB2lLY/F8OOO5CFkixLQ
Y7+LLkNOixWYuNuiQARzg+fXlsUseaU3Ra5TsVopY80RYIekqlTlgrP+Ngq7x8nI
NPs06p2ysS75yGL6pvhlI/ROv0kcyFyu9IOUX5YkPKE86jf270TifSolN/xyh7SN
GRcpUoTYHPlASUN9SVk0FhRw9k/w6Iz8d1TTbGOl0frbQbRfKOVPRcHpv1QQkp4E
vjDaddQpNkiSgwjtlCPtzZW06w8flY6F23SKGaIlnumZAMMLOawn8VxHbp7VnFEr
udGp5XR4ZLXtGTMHWB+y4XPz3oLIS57M2503uA7KJ3iZKgYiGWKL9tqBPDixMJxY
YL6n/gUObP+e+IeF/x+Zjq2vBgxu4EKazB3ezEFPpTRrPZAqQfpdw0BhrJoMYLxT
hJZbtV0jU1MI2d7GQDuhwSC54cIMMxUrZq4af57tBcrydSZbZN4J0Or1c4+LXHZf
efnF8214Cja1hpHpeuF/iqJfU3HwR/OUaYpCM7Oglx9tmmz4uQVQB6yy08yof2T0
HLvOqPGvP+4mcTw+tGoRU3uCPzY4DsiaBTle4lGFRL5H/qIlLqcbOK+gC8jsYIC4
2iV1Txwicqlgv4PEsXFEqzXH89vXZe1BdYR3pxPNZMeaPubFxUM6GRWWtHf3Zc65
pDup1wUSnwzK8PgetjcIV47C+AmVC/cXUcDYUWrDMPkjWZl0F7I6/8v2k5GHbV2x
31rO7FDIvGh9D+S5s2yrsTw/HckLvkI4/U4dimiY1Hya3oXA+PmzdYS5WWrbrKAH
s9wV31ZTRzDLteTHyD4nK0ejJ38Sgk1nCgQQIt0HRVPYtsi+ETa6yjnHRHSIgqwX
vqdSnbHqlXrPoBB5OQEGJ+GBMFw4J0bevFapy4sMF26m+XF5goT7qRWyxZKaZ8Gk
4R0JngTMvi9CsBqAAIKwJiEh8o0MGoqRUQs+IJ9SgRW4u3yY0d62bV5m1PiEJUd/
vaDT6RQ8N0cda+BILMIG1jL2CclKnkFl8J+9OgWVrAuDIJpUxQc/XiKcHmoTvsBA
CZLZC46+MYYlTIQ7rjuC1+kqVMeHw4loPC8e4oS3eanRerCHYKgmKAkbYsKUI7i5
S5cgwGw52F37BjXHWKFYfximQKV1h9MGIPLm02ZARy70frLAX8nwyDNSeReB5w5D
Vz8Vtlfl/UnB1gUejx8hWGS/CBOqDiirWkH4yNyqjmid54tXrApE5lo+MBTPPea5
AYrktL1BN+/4FjSxWUtJgNotNrzKIXmE/353cFJTrp1UPnh2DHRqrwcw4XrfstGu
90lSnE4HkKfxJZ8Y/o6IWxKmYzwcnnYZPAlE8ITAKAZTPhFIUQsYiJmPrtykxNXv
hfHLNLBCI0Umm3QHiTRuaOUx+jXGsbXHH2IbizPqX5iJRKdnLPpvwKPhDAmVKMN9
7XFk9qcfnUILNNS+0G6pplNwvYB5jCAE4M3XA6oVqR+xafdyTO5yvCPw776PS47o
ifzqd6JIlj8zfZUlE2DSdb3hqSgIPIjX0joi9t0PCDefDpz+9lHRTaImJWVeo+EB
1QMoyGvQgs4kPabPWCAolnyd3TVa3gIm7FOONCBN3B6AispTz4fydBIIr38IxISO
10MOBMnq+od0/OCoUZ6Rxl1QirmVMV7f+8XfScic3naUMqnh3VwSNL5Bbf035mb7
hjOi9BIjQuG0Dc0Rk0wgUpynpV5AfjtaSTPPca8VJOp187ib5lhah2c4OzAR5KI/
+yAUaRcQF9mcaVTc7c1sWXorBHALm3pg+4vgY6PXkz2zf+Qc40rM62r+OfVRidOA
U77Y8D+drngUHGfJ+nAj1OCLBVkepZoVR5HC6xscLtlMVR8AEiqmLrqR3b+WctEv
Lp6gvFUURY42pxs0ycwz8oizYi8SAMTxV7soK4JWB/jsaVpPjl5IOicACqAVoYJz
oomAbM9us+GecOiEsIFIBiU9LMwaN15S2IHpkrbf+maITNySpraz/+kz+cQzZLNI
0oDaUPlgPaHWDKoDlkRT7crv0Fzq0tICB9KIcT+pdTR38KQ6FET0pdkHn5C77Vgw
X68/rX5B34UE83Mwp4DWmzOCdMTPNQWVrtxdgVqJ1T8LYXOUCWe2Ynj6mhDVN6hF
VJFxP85nkElnjzem5IrSEx0duP6/br9HJjBnQEWQTPw0A/udSejPIsKsmXef5piQ
iVm57BmPMBlvnZFtCymp9BI1guot2LkXkO5kG1uPoygLy1sWuFvXEbnDvflsgT/I
ByMjVYJG2BCd+wK2FLLjnFHsh5MXYt100xG5ylzM16C/nkFzVj1dQ+/xiwgb2ReM
qb+zJs3ZgsyGcv5xC1ChoZxSFssfrX9ZtUtpo1ClzCfH6fUwMQDRK5VqGaNIymxN
Da6ncMz5o7sTVEf6bHJOPHQVmy/n9rl/rZHVUnCXS8lC3Bha+7ZZBJLl1Q7d6S4N
DTT2b4G9OQB63fsNw1CxfrLqUL5O28SHfaR7JdNOF4jVl5jxvHMmoB5VzEAWsmT4
mgI4Y3BWdfUQHUcJ1YjrURTyyRFog97E7tfjZp/Vd0nyJ135k77/6hKF0odYwwhg
k4XqiQ6hTAB8GfILKY0vqPmGiI5RHR9nfaG85dhx2FgUnGhvP5HRoY9M/BJxn3Yn
2f11uaUTdCVDRyRcDYgVU3asl5pNrbJkvLF25SRy0wkdjN0upBWRovGsxYXjPmwX
oeKrwiBuycQ8Mgvz8tTWxDoBeGjpXTn//eGxPl1KfGvDrmyuOcR8ekpPFyHGVA9X
Z7s588iIvqa5o/MuMHpSDR9uID9jgeYiYwd5jUj30QaqFYXu+Oh6v6noTfPu4a5t
Iw7FYJjKOfabzg3Ojmyd6xeIFMttMQs5ixdE2d6HHdHfBHKTVL7wPeYT7WZJ0q6h
l06gW/f0fkMBMti09A/9+Fa30sPtsFdz+j5knwcVoS1qFjjzha2tk0JQwk0EpJn0
XCZF70P6Wvbu9qjIY+jrcfUbPkm+Fc3DI9p8fZzqY19zLsM9/uEiwpOIp34n+n7p
VN2cSH6oYcXw0dza/2zjOcnyOagSPjyYon4TbP3mI5uWEDF8mtp0tZgy+fx6aJQC
45VzsuP+Of3zy1yxkmFAkz0xcI/Vq0Cr/YAUVh7UXNV5dx9Y4TJMFeMa5J/AHIf1
Cy2jvJ2l0tRgS9PHxgB+0FlS0C2BhwYG5eqIberXapCtf+1WXaEmVBVBqRQNFUEi
1zvMJOrGoOn+Ypd716lZrxzvHEmsBQV0URwSlNP4KnArnbyjt31wFoU1dB1U8neQ
TfKlXcnueMCI0xcrjoON49jgwgBP4Eo2BseHAevRh+itszDbgauS96puZPVGfiaR
9CL3KdHa7VmxRVhw02bHzr9ShsCkz/lRbXHD24QlCoi7DIW6pZyKhpBKYzOOB/x2
sWNLXOcOgJIDkMzfHV9pRTsdHHjtggdX/3TlBiqXJAAG5J8fWATmblt5MlCblPll
w6RjsTf1ePRNsOcTfyxEpOvT7p0Op11NjTtK8KzUrarRXDf1FTtLeWZ/FkJwSDQL
FbFEtmb9MjjeJkhoioI0DAEcBR/TuUqclFxDoWoJMNh+RuLxm8y1d2Vw6Ty+B7Ft
KRNbewIxIRAo8TQu1HtM+BaKxKxA2nITBZK2hNuDOKfUhD0VJlLorhVpf9cJZFYg
u3BCVifZiJLMQWPwx3QtRQcVML11ss42YFYRM67kQkqSaEtKm2g0A6s9w7RSGkJ9
/ZyUxYdiaLUoxXnpuTScmVa7SKWRIkctfUb9bO2+f7UXa4LKA1Y+cvlOP+ZjbZkv
I1zPCREBdcPG4jYHfirHmAx+SjurdAI/NGPjRX2VaFehb3FmlFQHrSmnwYlTbUM4
9rM1uTBpLZy+EaIuVzlCYNFFyl55+ETsFTW98gkQUaXHoR7V9AGokq2vmoAdoZCU
N8wi6QfOj7TkEmeYWYCZygqO5FnAhw2JgFNRCc2xC+f3CiKpG7mB9YbX9PCWpwXM
/diu36LeeIWJkDYi45M7qHsIYoXmcIr3eI1CGB9BH/BO2Sr/T+b0dPEsRuI0tpIG
hUn+CEOGA+7+4Hrf4hHb+ufd7YDW/L9rpUqD0U+e3/JdOU4U5fUPfJRGNOHv+QsK
O0qF8Sesghp+sd0s8SS4YofeTdVk8ufHlDhmSUfXaIKXsHkXLZ7Xsg+KF9IkTF2i
IGTfMz7v3ip452Eekw9y47JyByaQTZpc22K/iHdEhNd1OXqpKb5nJKdFELgupA7y
+e6JIJTwn2jE7fSVrlcCutaGAu/teVv+fadg1kH/rb8eGp9ZZWI0og5J6G7e9q19
BrJjM6dxYsP9J0LIlMTXXyblxGUwenFOO0e2UObJRhLegxcZjI9KAsWXTT6KpnsR
O9Kw/oayzncSOMiUBr44XXhhHpDWiswbDJLpTk13qE3lWgUPo1hzQ7ZDBF8IMGDT
ixeb5JPTxisGE39AybNTBRF1FC05oEazBKskhh4xxRlkRvILgeyBEU5CvHoJtHCi
yc4rikqHQz9Bep1EG2zXIFc4w6C6WNF1Vg5tIOaliib4BdF3wtzuKI2ICfw9hSQV
68wXPRK8GmJ9O5dWR5V1ceRPJcbWwZkDw1XokjjWnsrQ0L8DHAZ3z8776NCK/HY1
vG0XtpEH6D/HM4NIbD+QJF4GRi/3Zx5uh36ku1GAc7ms/45490pcYbtkJIvpvnci
iW7waTPs+AuhgF1tCOcJiBdJoQSg+TlaDe5T7ew/yNHybw7ejKPwX5eEJclTZvjs
h7HzQr2tpLH7J6mC7QW5rVsvzL5uiDFvK/Kz61ZWFwnoO5Ii6WWiUFjshn/2GIKz
Fg1/TwSC4ojomefcsXNCHKQVt2AlFJ2Y7UAKzuONj6C5qaZUfGbGOy9ox8REM1JL
SsnJXwlSogw1raYOR3zpN4dsShHfzKceyU12CSxsH8nRoQC6IwVCBssGcK8Fs8Sg
lf35y9b9lCfr9Y63UdP6X7n8irwv4EP9c8MGwZ8NUxcwlO18spr+advqqx2mu0wO
+OkmJKfFvBcorLyGJWgLOcXrBaaFwudmcUfXvlVxIBZZk/RMYNh07rENBcDVXnXv
MDEThTReRyZDAoanGZ56EuowUbexRG0od0LzsI2nXoxeKq19VTJlbGJmjpnXv4Ba
DPdkj0gtJhcz9c72uZWkdSgEEoj69GTXx/twg11R0d9nQBU7KHM85okVNHxectzB
LvKq8jPHa+3Be+GG1Ol1lKpo5gdLSyurABEavYHfK2ph4uWERoExGVIX/0UZcYLw
WUTInVjxWBGAp0DPIQ2pptM3nX54WfC5OMLjshcFISi80hG03pFDX+ZWr3m3cu9H
t6onaORKGgBZi1ANqk8D/hNdNL3r0VkNBObwBoozkINexxX2eVb2Vep6ZgGNdkZN
XFWqz473ohBw0VL0GHOGE10MR4vKo7tL43dSOC9HPKV6wmauYUQnxfBKT/SvsX3j
7xpeR6jVauSvEqbJX4tX33Mzrb4b5V+o4xgVO6DR1cOUVm+EEqlEJPaFy1tfJYHN
sytBG5amDPvBhfdvhH4DrL0jSBp9E6je2sApG/uYuu4CwBgxqpKRx2FnmtMkJXj/
NMWjE+xYNIlSU7IQcEAPk13u/E/hY3dqiQRcD6O0fpskjShG7r5mQb2cjZ1BjPdE
KI4VZe1GM4z/8qyxC0wpzmRztjRo7UFQWz6J4NgxMOs9ZezaZNTFzpxV07GzgouQ
JfVmq2pc/LcM2K4BYeE20jJgr8fTnwlMfcm0NDhs4wtnqBmVKk4vi5oB+44EQOda
sRQnJlK/FPWGACwhI3D2KerNPOcxe/FZgU2FFOeQsVL5uY8Zktb25xR1kqW932sX
Ex+L5XiLM956VoLG4LwNqYYgigWHbM+Hq/rnFrCNy0QC3OAt9e5lXiZavCIxN2yX
10VmPSWA5SRq8+tn8wWoHaparQRe0zruOvzCEnoA9RyxgyG2OCul3xtiI1k7ZarN
GcelpE7awpkZhIv2HpxsIRoOzyp2+qRIimtSsb/9xaIRmxZPBS31d7hPTU4zUwRk
GK1iLZBvUbAtkCoOx7wkMtyTyHUGcyzykJF0phD5wwwDXW9cF64h5HbHY1zK+865
x1+V90EKkDpB2pvjxwyf221oN6oX9kKsaIgEDY8qVULA+jNbrtU+OxEm7OXhRscd
yPNXkEwmEk8K73CaetjMyPWNt8d4p2Rmo5HRHGHh59/cTGrDqdbZ3joBlXda5T6L
dPaJYf0C9ikyzfzjsrMRCsTBH37dvGdR2GxA0IM/ckA6rtUtLibjBnFgsAGWrBDK
yEDjun/tm9a+eLZ4LvqvZbvVUqd8x7YO6B0GaIvA76i9iYAc2zPMV39gESC6u0Hg
T7J5pIQLQ/lNASt3j7/+VJ028uoSZdjaQYKyNSq2661K/DGU7+Z/yiytohhexq6M
uw9eXY/LhCkS1HThWvYJ8/C/2WHN2rA+lyambrahpFXI03BpnNImHUyOifM9jVzp
9T6Xs5s5ROb6UeWNA+TELr2amWYdvxCwu6CK8nKmX3Z3A0WxRpUOnf23juLBdq5u
TnsT0+Hvo2NF1prr201Mq63nIrx/2hOAs7FQ5k8815Q8iygwlIMXTjZjbSt9mjrO
rwU5Jsd/tLc/u4jBT2fDKdDahtfSHH5NdlZ8ym9a2huBmCOBQSzb503dVdxZe1+x
Ixtvx/0tAw3A7qq0xGZagyRNXNh62ojLHRvs2xE/IpDwTPMTzRchKFAmB8q4eXLM
qRY4FOaPopFR8zlqoSWD4mFHQoGFC1WZPLoAyUv8pLIlJJNDEVFhVlF7QO3j7Azq
Pt04n8Ib0mRAX3Pe42tEvrZPiJBZSMYxIcDz5ZqE0qDd0dcQXqnzeCH89TwgFizc
sge5UAJHTVjE99YJQKBClzEztylzEGG4JkdZiDVEuRnBSk5CZIy9WrUPmTaP4qvx
hgH6oSlIXwmWblrNc1pAhqXDBMPE9f2O6bz8ZI6yrmNxdeYF+tPCXFDn+yCZpASi
YbjRaH2UQPfDibj3DNyAENuD6C7vp2gK7clkzEqY4iiLr33S+sgsPNYAJ1NCkMFD
R8pjY2dbIVrg9bjRYkd3juw2OCFm+gwy32K9XFjoME5j9sCeYifzOgY8Ywt6iKLb
KoKQ9MP64fO3JKhLVAc2vwvUTMQsAPGZQnrxHsQlLMedxjBgKjm0zhjaQWo3BwZk
QGkmYWJHqo2BtPz9a92m6gDPbXVkqsmMQz8BQQI+slSFiGCqTJBW+NRD8+gETfp4
iDdbnjUwEn/MK/tj0zKqPeupMchT/0TggnakTekyJlXjuLuMb4XaSBWMjAfNMgj/
kYPxWMKrjmmb2HGSyF5KYMAoW7iE3IaWcKJseSvHV2VphJoBAC6/Tqw0/pJP4Gzo
u8EzCKR6DqopPuoLq/OQa+/MtwnO2SwSYTIXNI5plYR73/NM703kLlOH/Ipj09xQ
VhkJvyyjky5z0UAJP79KCfVoXC0RFa8nyD5I90q2krdrFDyTqB0Y9Qmqopo+m8ES
tCX3KASYNoiirHZg1IgrwASbnO4u0eO6BCwFmz0vaY+/pPDk01VWjLRG2gQXI/7b
veTXbrSDXIAT5PugGIRlETiMGPST1Oow0JLEElwO1yYFDsLtsK9PEawFo0lEPy9V
sVm1PbqQp502KnkMc4N4YUr/JW1Pccm+YNS3TUzGEnVrbP2dhyCFdNeMW5Zwz/To
nPgKPsL/tin1WS42f/iG4Poq2Wt8dinPxJmt0N1N/XNu2BH/+Td8xlwtjkMCCjIq
ybvkWDRG8qcjMneLcZxnDG9pUd3jWeylcYCXODzrzfZHyebWxqyvunTrmXZmv9up
MzYR1HTj+fpm0O957mYnDCLVdyU94ZQcJhhvlPHgRlmkGsnQAzD/GRB07LQNFSdN
1DN53uK9srXjEt0O/Q6159L97dMpRE1iJ3s4tbDSPkVedQF4zhOcKdqUS5DA6svS
aX4V1DBKCeBPsev3dAFu/qcRZ/RQ1Rpgg/Bx5Tw9PTXjhaYR4MF515OooLoGefpH
zfUcd50NoSZytHmVXAjwwSSoAU90euONBB4cJtKl5l0unW29ybyGaCx23slfXoad
u1+RjccrsXPk87Xu1bDjcNRPEMWUDvQXd6d3W3+UYRq8Oz2FNlFSrY1dePBU8Xd4
kze+n6rq65enrZrGeGAMKeKnW7iAoRYuQn2Lhb+dco3ajyq8rvvHdbyyWsQJGFL0
SCqqciM6vd2Yn2x1IWmRp7rs9RiA6Ysh6J0WVc2VvnJgz9X+/QatExC93W2u7fsu
upxQqviPg7KyJSbXS+UkqWHt3xTN6PxZF2202S0J+67hs9yRn9I5Jkblcgx1ikvX
B4NEDH0jAdakrnqzIPNRa0gaIfRlcXtGdMMwfY3g7iG6UwUpxhT6T58DYaqxarFQ
h9tWC1wKZ4RadxhNYLbno0e6LFTv7oEYDwMY5HiqQJ4h/8OkfkMG6mRI7RzcW3dO
SeoMh7M9APa5W9HhJu44pVFc6zPnQxjlfApPr0Z7dPJwMxHNVNnzW0PSf4bVjWno
8uzc5CjwTNTdsHjajTsfDVMEAV+iMbqXlz5/qYeI2dbSKCSB7W2J9/D4DI9D3klV
vQodMk/nlEHs42KY0sr/nxRhizb31lv6rhw83j5uRy7f6YVe+DzYHvn0hH4p2VQN
8rRbY+wipVK9iUuHD8ZxxQATd2DnF4iVVuCFK2VlYeTXVZvHNKB51DAPPyI1NNyl
WLCPlolZONQIXlWE7UzAqNUPZqAh+gC/870tYW6qxPxgU4qWuRXLMq4dR9oP33/3
jzpi54fgR6x9HJk/9N9Qigx9H8LV2cwBqTifSGmVl3tQ2a3T/0dHgeqltjbnPQpd
xSOreYyvH340OnSDSGYqGr+qsUVfUWF5AfUwa85O8zwOJ87NHXUqMlJLBLYKxy8g
atZAcD+CPbKnxqiWCtQvmKvg4A/5H86NhTqjZcAYKjBKRVMPVMfjdkQT4C82mmbA
j/6vhiOi7kfcgsBLNhPrv2Q1csIh4tv3MzGOqq5mnN7k/9AUMOMwnWlz4N17p/HJ
9fGC0USrdpvLx32ZzdO+2tyCEoswbZQmRNBpwpBseIldGm+u8jUO8VHrLA6YZUw+
ZhhAa84kABoQzTYvRE24dQpyhfu82mmd0SUE/uUsxEn1ZBOfrFaUNe/GDDF2Vklg
SaD3OoXoYjiXiCmk4qsNjbA6KJFZu65Y78+rCOSiVI+2x646cN6mQcHWIwlz1pnh
1zDcjvySqqUr6Vk1mRIqiY8sWEL6MDY9cDgxXCe/z1uumacPLbwF0z0g8xbqPQSu
mIXV4HSqWUXTZ970nKe96Mg6HCu1KeiMB4NfsxIeFyOqN81Tqfa4LBrUXAjcTcdT
pALLZFCtR9IgyTruXdxkccJmi0DdYZQf77q37DAXjJyxOeZdgz5MCmLlsnjnMgMk
EqCPzQmtrihbeKvaP9mQnmAeoqj9t8CYdRaXp5hPROLeiUwjlDS3hC0nJTpLJX3R
laCe+H1MQ/Qrp6ZNQiS6RbaJuSKUhVYHJU9JeVyX+lMCjiTLtwrFovw3qTsA2Sqi
yqlGSv7KWehDz0orHWnuaYixwJWnZmlFRRT/klBZTxzlZ6dTEcQee4v2yAAsrVWB
gBT2AW0NtDNpI9ywBR720s+GJ6Z3vG4TbxRjAUHBLQDDr3671SzfnSa6kUWaU5dT
sHIJ+E7SSVlgyb3sK5NnFMOeD6e4vN/ioNUVCtCyCNJ2ku2w8Ge7MJs/dNXNU2Jg
/DGETDWka2fcG5g0K2NZpG4FRFJb4L9edbc6lJ6pGU52MT//3c0bI+43TFLjFU3+
OedB58ZEOZtnKqc9r+873ela/z5CNPIkzIiZR/+kjy2nIQ3I6GuWVYoBDLgACap+
7znYDWKcXZ6z9702ixfAuDY7j9guYI38V5D4LFauau/l7MhZNUFBJ8RZh38lpsgE
RJXebrN5snnL/un7g0Q+Jqocje68bozBA+u3pzrR+mmtXMpT8GlGfrSl4RuI1ySK
gCsigbWEbhXm/RKYMRP0ApPyJR564IH8aGDDCNS84XFdTABHYHkC6xjqZvY4a6Bn
jk/jhm/yv0WjtyV2ggJ8LC/5ihpnFsQInGJUB5S3DD1p+Q0MVeLuWOtsQ5YF3PUA
Re5KC2vsTTqi7EObgE8OKRnb9KEQkYrNGbjLPcRcnF+LIhzsH4tIlUk/V5ueicAR
1QHJQWHfbIFIEPid/LGSZhvrIGCuQshxuDu+FCxgJ+ziHp6ApztQfp9/Opv5ynKb
TNvneVbuUJRG5xnZGgjBmtw8KebddTtqZB4gXfns6K+h3t7r10iIiq1pFYFuO1Oy
ZeNWSDQsobfPE10k7Iyy9ygLfRcIhg7O9TjWnPtIX+PmcJJE4e9kS4m+LhHxumYJ
t1ySvCCPWLSOvFiqHUxzuJdF4u8tiAsH9aPFRslXk1zvEUp/nVQ+i0R8QLpF+7+o
dyi9zkglLaq1cir/zaG/278WCmy8BdKKjAx8r6LNBAemQRA78HK8ChshzFNZuS/q
h+r0F219GONu3AdiCa5poNoUhCtB37o/tQIj5J4lBzdoKk1yqWzRC8bdR0tAdejd
cWnwmJ/eMNcG6iMR828kzhW9g52dY08coUsuk3XJ02wXRQD/28DbeH3EYBQkPMlz
2mKNqlw/02WYRdpPObR+V24NEy87o4QgsvAk6yA3W7m7dYncVjHwTCINkZbWJyx9
Ua84gRwjRxCBd8MxaWZ5+AurSael838EDj7rxLjUJAsLRmiNdY+LFHl9Sn52ZLyK
t4vKi81dfpdmuITVuVL18TKo3qd17GifMZE+Q2HXjWgltDfDmt+x56OrpthKss7L
QCPYp4RDHmxW5lmAFa7QBxSOL6tamUP2Z0B5ha7JMSb5fSob6F5GHWAjMXg1Vs2C
Y+P324oRev1vvAt1tLlz/eh13eC34hz/nuyUw7oJATjmqkGwtpsAcenT+Ae+JrdF
R5V88jNWeRhsZTb0ijkDYriduouK1ZTbIEkUM3XbAlTKwvXaMELqUYnSfHilHzgG
xxYp4AlhSAHEkHGQF46UJO6idwsrTca/mVJBZVar/qoppSVQD6PgDmM/eZjurxws
d2FWKNDRHlJlAsRfrut/DP4caZ4wVEegRvNcsZuZr6NJkhrOSpv0dIsOP2sRzva+
pVDIgN+F99rEO1/pMzsIW/5zgD4ELtio199W7uIgf8pLHgDZQdD20+TgifbK0bv4
hwAjlnXhYIzvc7hLHzrDCvXNFex9o5AxH1y/srP7Nsv7+j7OA7xC8LqQSeQ3db27
3nIbja6mJRsCmQPAURQh6spH4bcYP6u447sgbucg/MPI/tES9gzmHBHcMNDSo2B+
EAMDGXiosILhteq3EJMr5ZJzXgyfjzc4bpp8AU/4N7jdEkZwbxVXFlxP/+Z5zJzi
qOFm2oAutQ9VclP3vU8Rh6pWy72wcso4tx1YVN/qN5D7FOCSX1mh/dQjsAIQSLlD
pXHxcTvsTJ/pnSQqgn7toh5mKxVVM1HQIaDaoIBdiS2l0lUNqFTy3ysx0scGkjxE
BOjLpv0v1dvwVbqSYwGELiO07kfMYHbeSz3GmnnD2yI/KJ+aLWsO03c/Op3Zmmd1
ujt9u6LG66kWTSIFw0X3XIl8TeKySpridDXTAcLnpKlXBfg04ixmncsXRjmFNSdf
Enqh9Ny6/gpA8Rwh72+Zcs3S7htOgW/WWznW480sLlw6AGuq8FcVrsPHdrtLAqaw
A63jnsPO1osb+vMQg1Ja32c2bfMDkkhIhNZWK3dq0BHNPr/DssJGIKtWUQHW4pRy
iQOQg4DYwFE5DslVVy5vafKb562NbUk4rhXcaVWnwY50dgY2l5XVPxv7xXWK6vbG
MiTZ+z+dpdUUo7AAHS3GrwlVT9czXkahOB7aGF++qkI56JHApCCPebybr7VwvYNx
zPNKr6npZFJFYQrmePHxdp9ai5VTjMgq6Zd1O7RdnYbfCuWAL1WyFwS5AoZIgzyb
uD7VPrA9GPMHyKoIEsj6HuLhAAl/+yOTc/WzcTKOuSPXeM6r/ecKMYqL/HvXjfRU
C44+eeTvAMeghbglF8+A2lvneB26ZY7esBKlXR0/9/U5q90KONlu0rl0NddLNu1E
Nn517baqR6zhqpM+QV4fn630lFZ+YjbPG3LzieiWVfkrCl7HSL2zpFVoY12DUhAB
j/ay6cZ8mmH3GwDVWCEIX5idFrvSUT+VMoKH2aVhbnr5GrcGvjr3DEoEkU/YXG5G
kVn3uv8WNI+qiaq6sioMmvNYiVoB1RR1S+no+3vUf10+RVyKVpAzorUFq5ppZ8cD
eLyOqUx3XN8Uss/6G4Rm2OX5udQznE0T5Qo82HrOO5IILhu9XCpjUW7DtHaYv2z6
8hT2Mj83mK93h0b0IiJKAXKySgZtuq1B1J+ZfDBCcshWoJ1i7nrXnqeeDjdTN70e
FundgwjEsel/Sx08SSBGkLHENkcMo01th95lloBVWzGIV9XjYZjvbTS5CAovCiW2
ItDQKS1thaJx58hiMnN/ecvCkl3NQS4ghqE33dhr+sKbqInwXB3/0NBt2cs/+4j+
bZE0Im/mltCjmWLprVysHhpQJG5J2m/Cj6LJ0q8RWGmoikmHaxqw2QDeOwuG1mIs
caO7e1L5bZmovRjiagbuo8QcIQPP/CXOTFHPmDa0f4RIVoOLks0wK1kooMactvyn
Hmdrxl9NOu2UWfFyANZIzAngWpZusLoJptOyxTfb6YQKY6Fr9Xa9Pv7lMlaDfUBw
ruvuOlMdwaEiopsUNxRz6TOu5tLD2ug8oH6wgUrVkUZOdM+7MIT6N1ek03Ilirwr
+M1xkgQVgekEe6QE28vts1XaNgRXE1QwypTjd/300vmP3UXPpVbAQaStLHZjByQC
YBcSIF0/h5pGWgZOBJxIc73VB0SEUYoo7x5VAxD8tPaOrEtiPdD+1T4T/GLW+5J0
bDizvgTs/vrKUefll/tFpZCmV0ZsJobaeml//ZfGEOMbUa2UNGEfqf7dpCddFl+r
qqLNzBuML1zFcT/MboNdIxt78b4KD7fb5e7grlzB04Xmh/1dfWTPuec9M5cmGOZL
ZsCLZWaE2ydyTRNP4soVMN/Tfd+RPN93aznzYgS6rmiWejjY70DMI8qZtCw/8CFe
o8TOfCLXuhe9t5iXBv0M/JMbuPGkgRsj2H12p1Cg3Nj8plwrZcMWcCq137NLpCSK
UfbgVXs3lgIo2wDgburUiG/ccD3jTfy5/qmHIaGSEQIbnBb75zCz9us7TyS6IDm/
2eiJxRIQT0QytinnQmvLB729WYmF7q6JGqgyHHJ3EenylmicK58ZkmvCUpBJEQxe
OhGbUWj0+NS8B1Bzk7DzZSuXr/CYVm99vhK9a7VHd91lTv4G+LKRFGwcaKZzxxrV
rOMMnt88X73KFn8Y82Znf4L/9jjAMIX1pV7jorojHjCfXGtPV307gezu+8Fmdns5
taHOujKi+FQhgboUNwlrALkw835aJjDXGigAGN9nkDCTTc3MXW9HTNIHRQRnyyqY
2iCJ4AqZRGcKbfVScsIUyCzwkDqb7KdJtzGEyWw7DqEXTTCStn/LCUmGWCyQEp7G
e9grptCGAhAiAkKZiCqpbjzIzZAQABHmfsyXrVRE0blipS68xbdBMK7Mc+4q9s0W
9vcUWABn0PSLjjLidniCS7rmNQdEuxQOvAr3gkAqovRo6L1k+euTO8KZjIJtIpdq
nuLSlj5w8UOE8T0+TCoeni3sgKiCtJi4C3ZUqjTA5h9xz1Uggx06iuLb5TujFbWA
l6o4bCVClOHnotKRYuZn36C6+UKhbIBvqpUWA+vtYA7ArOvKhGynzZKCnqRbdE7n
vAVDw3dMPV9U7g3mobdDIbKU/4aAQ2H1CkC1kwawHItPlEDjNf3qCFXPegnmt4l0
APTtV4ItW8SLVcXaxcJ+1zbXuOxuHFQLbH6+UoV4kmKz83R+DRzLXROo5PolUbRD
NkWHdRETI5joxqrl3MOHrFbfWyHuUS0BubcVNmyN6cjh0C3HzhlGsLp6kfftJQ3B
bTf10HXjb6HeEU8bqcLfFwpd3yZi0BK0NGvch2OHcXD0IS+gpGJUzcCFcIo3Hp3X
oXbQKUW/Hkc8VM2Uzda7TTWPMK4ZPNOLwUS6ykgPY/RvoVsS8VKEJKVzvnDCYsmy
NbMVICfCh97WMaJBoZSfSNPANCga9QnJNnTTpyBxcko/NhSOD4CkArlZELoBI0kw
rBsXwyIt9tqwsOTLn9F3WbyFRSW3lGHxlhj8c4YI3uaH8odjcUTdd4a4M6T4Nor3
9xr4rPiJCoCNWSvjh5vvlPU2lSZZSs8tPeq9zYjDv9WJuWySlr7VxY6FSjFWAQjR
jSuYwmyWeKijcgetjKJwocLa6qN0Eb7YSpMkp11PAwkAqEH+rI5txidz1dNThdaW
8g0QTyeWhArwwkIN1Odhij8F7vti0Pga4f7K0/BRn09DjBNfpxdC44RXpyLjbIsw
qm3o5ZOLC8b3pWmQWPi+AZY/LMlJUotJwnCRmKs8l1RMGA/425+1Dc3qgH1G6++g
WFZblrO51Dc8O0fhvM5mfBhNaBp66XTmSCTKMW/53TnO8u5GPCEXJyYkOj7bGC+J
D4Yn7UU7HXNhNFau4kbhs2SiZjM7479POnO3KpQnFh93Zf+WweeUMrZs6zBH6aX5
4nmU3ozsgjR/lnZ/lErQS1uJNTy8APu4jm15abJgom1I4pKUm0i7SGJeILEv9YD6
FVHCfCC9+M1LRk8w7JMJF0d8FLOGHufxD4I4bolwy916AmHBI0U7w9ri9b3vT6lm
2yLhn2AsWOy1A9BxLtgRmSLMpUMQw1uRbhC7M5DjDMw3jseYIHtjuZDShBrPAToE
VlI3Up2Ro2Fy6L/+vMsNtFrvV42mVZjg//k7CCKpSUTYuIaUIOl8+dWS9cA0ZGvO
cQVGHiuT9y5ZlpJkKg+6MKvA6OtnbpfFfgVN41v6+hJpSs4v+7SX7VAydWGD83Lr
w6TVY1QlKpVE84x6Kv56NBQcywokN9brRL9OV6mATg65/rfim86wFFbVEYM8u6ss
BBjTADBiSoWyAziHU9NNjacWf0Bzh/eWlb04c/3fLMT5Bvl/u+ropIZWnESiuEP6
+0tvR/THWP0SP8f/hxPOzH/iJ7Z+NHoNCN8Sdjv0wVGMgQJ8BQRvTt8FMM7pwCbl
saF4TZbZ9uxxpV2L1/Pk6PZqP2+kCLkUGutEVh3YO44G9Ke9NGPb+n6Aj7pdWiNh
KMZXK5WyUp0/4Bcbggrzo8XOsWpSuVriwmgeohMs2ESUGDSTHgLa3Wx3SUaCVmj0
tmjCA3SZMtaYLO85bx/PDPA8tan77jsjMhJZq+rX9BaSKaTbt6IMakFQnoU5HwJ2
FWn8E+9HgoAdM8J0rLKtGQSZGbBZquk7roqLiDZPrhdkX0nW1+2A+vr5JO4LF9yy
cv8o0dB4ougQXt5dewdjPzhEFbVMsgJYTSLblchvU61Yxxr+qz8E94NLsTBy9dc4
criPaPQW3WegLzJLX80G8kHKo3p9f3Qx6GJbVMC9g//5MQLsnBMa0knns6dgm4uo
v7QwLhmDRMlgGwgYVtdlzoWvZTM3DjG3wGYyJx1u+XHr2c8E77tTPNWhP0qhcX8o
bjj32Xj9AIvF0x7VMqPMxXrFhpZQL/cpdnvKjvHz/KQWJ0oLDpdTg90DmiqBJJU5
k+UiMN1wTxN/QgWXcfkiRYT/InIvoZoo8qJSK1sloI+trGO5pc+3UuOhjI5rOViY
EqikCLxp+OUj/Eepacv+QhU5hC4PYNxEdyT1S1DwtVPO5OLjGsJZfiiiSrX0m92F
zmyaPVI0DtOFy9l+rO93xkC1IPFfkV/Z25dhfa4kMdZGXDyc5yOdOirUU0RpcG/X
w/Sa2fLG5vJwebM4s7N9yYOI9NdLhnZYVXz65IjK+tEY8z+FqKxq2Bzu4vArNq87
7EQZwCrle6U8p00NHQMxajvAw/fihvTj8vBkx4WOvO9qh/Nnro9EsfPLlgtHxzW1
J2ja6//VdkXVIzSSpcViHFEUXr5ttOoo6YlVUjNSaDeg9mxd6uNDKqhzVl10Mo6Y
LJvU90StSc+FeZXqPrCBbyuoc4yKnVojLTnJV/oeRl0LuylLu1uawVoglvWDUWzh
pB6bdZMTpOSrAsHdWwz/jm0zEVc20tBeh4IKjS1vrI6+zHI7H23uL8PiP3JyJmVB
AFi4Wn56uJmbjP7sLXGneTNUe6M0SS4vGfdOOI70OQXjTuwDET946UX/Gh5T6bza
5kiFIWH/HD8CIVK4rhQhHh3QxonG52DRH5RYtE3FHTS7oi6A2PXzPYbuKdrwWM1l
IrWH+tfzGBtGC9fLt4whDdVHZWkJxMC+5+BbIeFHd3t9BJCDAQjysp/NGsVJViDP
DLoajbUK4h1yuMrmt0tUJhtnr00B+LOd0D7x36ClkGa+ouQi+tZEwTqn/06BJ6GB
AXtKOm3+rE9wbMSBdR9aP2C8GfvolA/GkucZn/+FoR3QKsGCVBt2PyCgmYr7KBHd
X9wJqCtKWFNLCAR6axoqOaD9AXwpk8cQk4GLrnDgSD6LuD0032qr7poXW3RiADPt
0KmEEG9Ls4MiVtY3manpGJVsF7AXXr3l+tiJVTRaqt5aG6PpBs8+IYLrdvIo9mB/
rwMkGz+zyYBgkWP7AMuWpCE1EfQAeGMRLs5t00Oyke1TJfCYUds7KHnjT+SQqZbJ
qySq5eWhbLjy9EiWETOaN4mcbKOSdDBbm/eyrvEVrxjQ93RfVltPlpxdgWM2bhwy
6U+5aE0VKAv9zQZhiCH1ON4sX9CCH3J7a3eSb3xpSk32vJryt55BwnVmqt4Z7g5r
kHZbSndCc/TKQzM0e0PJiT31YjL+b5Phi52Sb/jQGr/0SprxNTFl1WA4x8HvvKLK
jOkX0ZY/r4MUVezDM3H+W2bPw6AA2egJjbKHSI1m31qKNa2xJE35up4sZp9h5gwq
aquQEJHZsPuF0H+awngUltJRhT/XmpeuIxAmC4hbPfDH9L5Mj6rcb+14GvXS5uuQ
JBGfTq7S1NQESBQP2VYCz/NUrOqjDOJYZfmK+3ECt3/lKXn8XKVntm8AljB/GPfu
V0sp1K5HEz48q0+HdQF+uQ8RYUzyUQSjgJuioO21TwImOAQ/V3ibL2aBPM66qfaG
7IdrCY71sUY5+Uwr/B9geu3j6+f9jbmNaxVvYCmwbCx4BwUgGO+6M3wGvuBEQspy
Ke9YjiNcUrBhxP4KplqbXuqWIkQWhqdDVus/SRdrqkWB/gzgHiPCt+MSJZOZnpVo
b9y0kAf5QvCrbtN38qAvpoSpSXUWJFl4dC9Hy3X48l6sfxYwoh/CYqea2tYppzmd
8ySEK9GfZ0YWrRjh0BhvLti52waK5KefbtgmeTawH2xva6v0SRlGRXogPll4YDmG
ivR/qPcSa8HL5gNm2UXJT8Xkfs7Ha+NJoqIN1o2Yi3+xAlpxIfI1ob5uebb7rwEj
OrJLVAjjpFFyyI0OVW1NmuUTmjyx4wrkf4HJVLREcnD3x0VSZEk6Q4e+ZicAK6BB
W6jPVlNqoqh6vxdDzP8hpoajSofiOnrbTqTZlo3etnycfvapTitwjwPCpiK3U8Z4
l6FlmOopkPBM6JKkFES49UwxZYKs8VN4+qa0FnJfzAkbv7Q6doy7uDWbqLlrzIij
LMkYcYxaP8TmTQ+a4rEjGncZ/tvhg6TfbUCa3AqMPpZ1K4JqlKx15BxTmQ+/U0qM
fsPdEqBZ4rqmrztVwXexTY7CASsLQRLiav6dOCjGpcw3xveG6V3LEu7c9e2ibpoE
Ys6Wj3tybgY1EEA+5VpdSxqzPd6YEFbd3EXaWffXlyfFwKM1R6YZqZ7Xaedx39oJ
BHhrz7TeBYtI4QfTfKl2LNMWtAfwnGYJcE7xgEZE1UrYK6B4NBbhUMnb542o5dAF
fV1Px54YO+R/d1pMzRc1QokxSz6VWZZQYM8n1EhF/3EM01poL685kO9RsyGXnCUz
iL1pdTNmY55qCa2aUoa2nvdUvOWN8a9FCknDJP7GfFabWmDxStrwjQNrk42J/j+u
ya6zS0ugCN39DdTbbA6vuoodIzv8YjAU+rBsl/JliTWWCB7TbrDDySru4nodAlyF
1wweeMVdokzlqC0DVzRY0lQ1b70jg5186+hbmfzbK8us3R2nbQKzBAS/0s06Nso/
zAFEHcc+z34b85etFCYtt6xd+/BO5hGEIiEq1MFKl3B+fE1NIeexdAl25G4Wi55r
5xXbd77BvHnNbfIdhzr5Qd9q8bVS9K4AIFruY3lqD7sKB2iaaQiim+gkJbHqJXnr
KQ9GTjRmWisqdZIPsPCTXrByeizGDo44SOfpU3orLll4+BrrBWWCyV8Zwr0ReIAN
N13TnvESE59ZFemhMimEgmOXE02727HOJ+/X875CKXMLTpAhHre44AyptdDZqaBi
cHF1A8uch5niKBZY63ftSQbjgqR31KXtEjITRyHy8B903ogQGEyCngdBM+/k+V2t
Piu9yY0UI0PpJovsYtjbkAmxfLt2sT/cHQo+YDX3t36b0aKggikt5fl9cRvutowe
viCcbxfbjra043FvV7m0SeHX2kEdNLb1XpXoSVVuqy3iJytK4lGfi2Pl2Wrepwa/
H7Rq3Fj8HE6HfFSubbMZIfJ6DJH0sJbXgKjHbmW2yDeyhyVOG3J+AZdygoMao/pe
gnJZEqItljLSyW/VjkF1avKDEQMqIm+zex9RSkdi6WIF40XypuxNEZ5H5/xsqhlY
+FOFYipbjISNPyay9dthl+Wqjp41PFQTWiLNMvbzuTJcMwALLBfniwsmB9wekRzV
iweifu5Ue6TgU1ejBvkKZWP0oFNFPZFP5SSkhx1Xp72D0iZGUvrDiSh/k4yyIOev
CIJwz3zK6+g9ADgYoRdZuwgVqvwHNCyG/4GTL0tv7YojNUmtmFKrY4t1ZQ5Xjzwd
ZPcXuW3n6GZMJWQSwp2CT5D0r5gANsg9j74i5RJ6L5Q/CT3nJM7NhztNSKJtB/cD
4Qpe3lSW/OwwTa6dTHpHCFWf6m87FMkVzdouE2CSpp5qpNXRXh5g+OddRKueHLKJ
DaAZsHZZUqsRnmsEAcOWQdXvn9ZJ1pyyNMjPwytypx4aUqbkUktmb3GGsNUPF822
poIDwIoPhJpGgoOA0EQwyVXTQmjJOjaC4DFS6/H9InyJw68IDjld6t55zs4Troic
iDuxT1fcRyNhyMLFt8/TE8sGvnbfbMnxbRHxVBN+DFqCixwIcx+deyfbYKTXLtH0
UU/ptUzUGBVrjfmK8/WCe3I0nR7TNUj5G3qCdNPxfIAm4WqB8YGrVt4xk8/ICWdf
tssC33Q8LHTLUIgidprfaQxkclRednG3xgEm5K+wnyn6umuYeLY8bgbQsPL43Bzl
cML+OVEXCNASkxR6WoVw/QBp+tB196u7cbrgvvZrIo7ezNnstlClqfBbZDn4df+b
GRqgHyfL4abiXkkLEEsCA9lBP12hamB9pZ2dFWxexxMUPXNxkZ+D37sNK8p4sCnu
h8pQ6sI0TZLGF2RGy5Tn/IURbOUpdBPpwa9O7kb/t9wsGMLcHjB9Wt+bSYfvJ0dh
YkRQQ9oUpj2+QjHf7wIlOZcAka2Lh4pXYp1GcF+2OG4zV/bU7uBo47EjciElYq7e
ulziLgdAEO9LkKMxSpgk9ASFU+sLkhbg0wvDqBYuCkGnH3u25UU/JqiiS/LQcnda
H885OcH9mTTFEmeyrLf1P18o8oCtTOAVQNVGE0EBMeY2+XDRQ9Gev2KI7+5T4/9V
GPjzxlda7uNHkhrQEObl/DgtUncjDxOrK72hkB4UmW/ATOrbxWZBagB23zZE/da7
U0p0WLo4OEZjXdOTP+nhEjQpmNan28nCyPZ6icbCH3gL4zZ+kX2gf6UJ3gyBvBIg
XsTLdeW7kAvknRDLsDOBfPdsD3OdTrYNtK8ImTAaY4wA+Pfzn5tXaZ7hlGikwVOa
G7+nP/PYBXhD7tTFV8aD/ARiJVi0vwhKIV1/mfE5lpEGzFvCQb/EKBYwXxQMpvf3
Qz1NXwdwPi6Ur4z+y895+CSeD5RQNAJGHAa98NrjrdVFU3J/uMpYJ6nTl1ReRQ75
7KewFJG+rfHBRace5xy7d0oWiJSc+D2fw8ygIZnFfYQAFykiIfpO1k999ya1sKRf
NPXzH5h1BzisUrSRawa9CLnigb6YO9KY7IFrEEU7oCm7YUONYbcDHOqQCSzWkXzh
90DJ6SCvvVPFQ4v09JydTsl/pdC21t8likjwis03/bajQ9jEws42xKb4F9ELeQId
X9FIVb7nW5YQjxSoQaJtjJoAQKY4l+bGNt/wIZDWuulrEFVx76vjA4cC01kK+uQV
ajBe+ZufYiD1Tgtc01FkgBrJAg9PN1jBMqwaqhgR4O+Xp3ebqkb4tbvG/5uSWEEJ
gXFT2bD8tHlNFn+tnSk2hkVmVkHdIcNguLK9HuWzoP75XjNeCGFb3Fg2nDgdk/MU
2aXhxVK3EA3G+sDDvKFse7Q5+2kN1CQWTupYpOq+NvER9bb8F5rD/B5cR78jIZVm
RTYuWH9a6c1EGE3dXEZNy3SFsuEinR4MMhMboWsU2IpXK7E/iT8llzyEv9RIEtV/
fM+3KX9Kh2rhOlMS/Rh8ljuuyx4Kyv1yDlIACHknRrgo+xnjvoR69cMsiKG+uxMO
3+TreKvVrcl+6J5DXVyEwJg2jmDLWEnM5+w1IjVOEfIvNmPP6yWmHrHwA2+VU/Ph
AydnFhfDU4odk1SUjvPJbxhpeXdmzVncMTrW6rs6KlgerwEHAEtsN+4XGE/++Y99
NVHGIYQnwYrf1kEKNp++e83Jq0LkQNpz/As9X3HWIgj975Kaw/mZYUavtHAS7dDI
tqk9fhR7hqffwICS3xdlzoPPqnE+2loiFPnlxSvPyI3X56h8qDA0KQpV3BuT3ESO
b/JfwFunmO+k7RsqzeM0p3sttk6jlYf+Zdwscyp7ZiJJU/1vpeH3S9KjiSiwSeew
WTV3PmY/xf8YkiqJ+2KkejvJGtjIOLotVJs0+w2G1xNsbelH004jpVavL+LkZTD6
h/oOIO0eAG/UTGhQgL0ZNAbP4sZZnLmG90t4A/N2z4UiBmpFW35m37N6aJpDVYxB
SxgxmAnHZ12FlHENaADCXcWHYEcCBKJ5xfu7UGMZJEKoJ1imdMSaE8LZ7Ud81IM8
2v+t0USLTi474l294IwMpwk/5QSnkI/CZziQj+jnxRXC91a6Em7E+qvVSG90Z9+4
w+wVpYEi/nqHXi2sV+HHJDmVqDTyv7ojf9T2/PyNT3McvMvAKzTviI9FdZ0NtBTh
PT9RXX6y4VUWKUa+qTX5rKeay9dDkITYMoxDcmTWKnWOTJhehpz6PmbdvzTNN5Fr
592qKDXJ27uhjBLwBcCYv/d0k7SkNpaHqh2JqO23Wy5YqOL+BIbpdu7EtJA2m5Kr
IXYV2d/a6TpG83m6yfZHLiLtpGDZ3i4EQQWf7XG9iHbj/fhS8mGaykS07sDWGhQ8
ns/k9F43dqU9GUyGeTaxkpFSlCzVPRijmIllz8emwEZMFB3aRT2s8wuZlIvLhaoJ
/+x/efKAs0xrdE+je4CSnz0tp78Ewvl2nfFlFCyZXVSWTNOiOjO4SHB6S1PSeOOf
MJe2QBMQ4Y1EJRrF86R/ChbIL8d6EcXC0SFzpZsTOw5I2rxKVG6YC+VUdZzBXSnf
96Gou2CoHbPbF54rd8FA+ZWyZjX8Xp5On3TKMnQRaFVBnG9Ifk8tOY/Mx0FLZL5v
mm+zdv9F69MzLPyU2nTuiUoZvX/xv1uVRzC9k7NrTsw6j8I2ewetbIwBMAd7195V
RYP80UElmmA6zNjpp0s9GUYyeSidrC2IBeePJ5gNAJ+bxCJPiQLtHnSejqLKeK/i
gTRYrJDGS4ax0B2pW1qmGxKcmnr1k5oiB/mc6LTYt+PYwaOyfO5rih5DPSb5Fxpx
b8KuecPYKdyp7rl/U5JIuOK5Rx9zBYbJCWS+DzhADFLrvBYnKC+eRToVVEy00A2Q
WwPsYT2VkEbSjwAPwqOzQd9Rcwp/rMy4V4Aps8k/zVjkAtWQoZIWQXeL6q/h3V4d
GUHfUlKn2ABf7UZyz7wAHQJDToJ5S/liBmXldzQ2fEVKmr+yXyANsuj2B8LTZ/b5
FBZiUYONXUjtRbHq7n8XDbeSor7vXGn+jQNafFOpHhzooXUlnEiY1pG0tV3iuQBy
jIxklXE2JwuC0wzrNOyubBQA3ojTrkTDt8jPl4Ywb90C5HyIun8XmEsCcD9j8Yj4
L9dTHCc/7pvl2VPfJ0R2+UgJYxn5DtEuJcqfu8wj7QRzkleO0kyxRK6b8tnauGM3
o3GZIZTGXXSybnCprVdrejrWm6C6/E7b4Pak+C8EdJ2RgBrETA6eMECqpROnDHb+
rn0jlVMfo+ILykk6nPuod4090BeFNFr8z8fhbRnAAEq0grhc6VJ6188FI/kSOqKD
dwCRxVBl9xnUDf82FCdEet488ESua9PAae5F0bRdrK8Wh86Nw6Er3wQJgdBAQxa+
zvJt0Xq1SIh12HgQztz3Qs+GLeOpFEpW3DccLXxpkU2eQqxGXO5O+Bzj4NWpQlqF
zsDux7tH9l2q8zVZKTKsBYc/eFYuCpMdDNJUt/kzH9ZyCqyTnznyleCT4dmUe0a3
VqX8BjV4IpN8LDab8Drpj+OC6V1zPb1D9/ODRzYRoj3rnUdYFU5We7ej+qRCe39Q
X5/CA03ZFwZrLuD3zNBUaW/uhNoKLowwHlxXSIrxlM8Zq00DLgoklAmfJWrKsxnx
RijhK0vbtC3oDiZKx2rb9pCNsU/hss5bX3N720C7rs7I14cSrDDHxnZbCKES8hI8
OVIIfGCUjHjxdBwAKMR+Uko9fkJrxG8CGFg9by4PAmnVKX5OQLWp/B3iInZJ+ekr
bRYJlHqN0AqMhMWCgPgXwvqZafpC5RDM48A6qZzBe42qg1XYGnD4C2Gwtk2qv5or
8nr95/ACKX6DrMV2gcHpUab9RTfrwoArJqqMQ3P5EMV7YIGRnIyt8dmQkrbPB9x8
VNJrT/B2l7a/S4jNhegOColWa0TnnVJMunC7UmTkBFLEybfHfkXrUL6asbE4bzFk
eOsz61EskB6f/3qkv04FAHH9BJzUg0qzwZBEGH4vrTHHfrwQeey/afTMa+s4zBMc
1qOXetavK+ZyAGx4RmMJRs3y6BwzH04snu7phYto5c8ilgfkfcpMbwARJReHHrxN
eBOSXLqX/fRfUJDo1pgYWrA1Mty1DMDVy5KaCy+kdRxaEoIOyywTWTTa8sTVprUO
O7thGLzZTIPxqFSWTRVKTnozDLxUxjG8R4286D0TKxh/+PsOgNCn/oxT8bm+ZQIf
N2Nn61EkabOLscpa4rWtj7wg1nMNc6CuyWJkjv4Vxsl8NwH6dqKtFr6xJkDwUCR4
kYTqs9esf96WcJl4X4uhP6RP4y/pDZv52NjitK/1Jg7DTalMK/E1SPxM1MO38wvG
Ivg8nyVcdNxluiesICyq6dDzCjdxLhyu7Ji00CkIAajUItTHBI8w/Jqaiy/997jx
nxsJHKps1VogqkADPzEb0UWPITBbZe5XJFRk9jYEpHa+evHZ/SYwfwyqRITWQr2T
xURMexyltMVwt9GrELNc6mptPj38iVUiq7D4nJ2Z63/5BZLNjBeEGfcI2wmgXCqW
1i248PK88DaLgOini/QnM1PcDVNi8yV0WHqk2kkcFD1pJNNzlzFTv/y8D69e2HCq
NGigcYPU9r3ZM0gu4zno7GTE/aV32CXg80b4IjjnI6Cmu9vNQWJxtRw7AvMxf83t
moDgFkGpfdUa1tqhzCIv9WbMnkdxtgfAaWdnTVr15dnxgT7yUrcEbhRbajFHh2mw
0+wR9nAuvloiiYUl57k8Xlii9QfJZ8tLLvdlU0eb+twM8fK6WchddTSUcn48jGx7
+yANjf5QZRg1lpIfPaV8loEzNzAAhChl+ihD2RTIiybBiYFH9NEbiVrxyACgyqZe
iiMNy4nydk1yG1vacRobZ0RElNIh0N7Ri06gLVs1HJn94osMlQ22g69ndBeMQgT5
OasXIJrXyncQQVS89V7GRlR8o5JF1YBjzueNZCP6CA943v3Z8smo+dks9NLME1en
Wqyv1/399Jc2/Q0QBz/udtVG9NzOPmVunECH71k1+wWPNQjOAJ6VoTCbq0ZRThuH
Qi+U8cvTXa8mem7tbkdgi85JbzWabpnMtB/C4XCA8QIkU0Ekg5n+RxnDnSbfpQdA
qlhpADQXQATO84I/EVOKsNHLuF4YHNMNbs3eUJ0WIzJhhc5IsWtK2RweT4Q+paOX
50Kv/VZRLi2BCRNEMmK1RXUJg9MOwzTNJu5hWcpcA744KRGSytQ6paf4/uye3dsp
lvPAWgpwK/Nu5/BiOSaRctk3EDwEInC4rm4Ok0uEg1tkQhrtCr8rMA/M31iywYPq
1qcicmQXHQkHeF4qEXeBKxKwrpzLUlTS2CjQeHp6d2FYebikivuI7Y9HUVxPVEDK
Ph5qKOAvPFsRWlE3fiNYDjRPaFf6u6+ALPtzIRqDOzxCghHNMYAmWM/5QRuu4Np1
GMDUxjnHXlJhm5xOlkRD2u7e7T9rmJ+SM7Q/xCUmPTOxYColg1Ck5GZM529GhryX
AJiE+fwxN/omDhGHohl/CsV+MhysbxMVM+k9L1U9GMv+pXw63VgCZJQN+HIWpy/F
9A+KCeXijxIRIrbudvP3MaI9b1AIp03S/zj8ZDP2Cg4fHPs4YOMYTgqzUNrSl+BS
sNGSsBqeR4bTTYfHbxD6ZfLXN4ZZ8tVMik0eKuz6kxWe7ea0lh01y9vmjm15lnV9
TBh4TrEZbHqkbvUXVPt1QGiExpS0Z/HaqkIUBn/ykbLu7JNcgzKoz71QGL/iHHUv
KmvEXeFxHKs0rKQ6/NRrJXEORC3BQP+kAhK74+ebGkJb2BNR358m+KLQbNIrFjEx
eYGBKiE4nsFAS/eQiFAfxHL1Q4njy85ryrSC/ODn8TF8Sg8+ndyBiHCGM9cTq5/y
bKVeXmcj2ooXb28vefF+1BT4rBXWU2SnRa2Q5b1/QLJMEl+jqWVkuKr+75w6XoFz
w9maTJNoxgpgn3xHLODSY8qb5iwrXKcpxTa0FfPpt3mxRIMiE/htywXFvRkhIiO/
ppPIIQmPK9/3xLmYRSR8W/wNSS4m2SoFnBY16OWJRQuJ0+kPzfQsVGKv7d47O+Sk
QPxLgvS3snN3MmPqcFsuWAIdfRInldKhX0+3XWJc4CZKC0ybcS5ZkwBAm4l02Kpj
dd18aZm4W58zS6VkpwjpfIbzidBLng2dW14chS5xZTnCISEuHh8WuclGWAzj5YFI
Le3mUqVcGj/EElyyIAKKaO708eDK+N/39LpE4vF+Gp0XGIILayjXvGt5KxCSSI9s
eyMPnYeF207vFv9fpIDYty8dwF23Y1b1NGDAUgKHRmYsNhYyyfHaR67TycmDpZwh
4dla7fKNAoC4BCdI4iPbEL7rjJVMFCohBzNnvSdxiTnGzQ3vAvLJHEjxtOA/6B67
P50A1Gx34SGIfiRGeiLo6kkJbsypnJnwK1MKMDUjwP0oCmTEzZ6nPEggpd/GIJ2H
FL28j0WAr/HmCwEZWpqmc/1RDVImT97t5IZu7ZIT3eaRo4W4GubylSyrWluHOsL+
2DVo4wVLFZVkV9QUBc9HCLsv3d2bPuEm3JstluMZVVR7PWg4AtNy6ntWAOuTfElv
JBW4NUPZWEg4DddReECYq0dcCw/HJ6A/fj77Lb1rG5km3v3Q+l5vCxz44MAUfqNa
MT0rJfJrnYJfvTDhmdv6cXrKlmGUHYaytw4BEg8LiGqVkMFMfc/ZB8iPp++xUbje
251SLe+cjfeOJDzsjNvWvOiOLNPrq8x7FUAzieShlwPcCpcRnO+4li/tyIwdMBDk
PQ43HIf7bu1u5TF596D3Bx1ksgcqulsWxpfFXe+tPKo9FWuuvsL3f5G4snxGfBEF
cSBe8Eau6H4zMFU6rI4A0ti1nsqxiQESYej4lUD0tcPifKlZqKPK5525fHh0OH+p
CJCyG2RLF5r6nTza6lpg1ONXBSz6He21DWQpTChvvLb7qGeKm5qVzNK/p2zOPexk
YH/tBQH0ioVF+Qgm/mIYYt1Gm0mIGx8V1furGEonoiZYgBwOa7MzfRLofhcetUVS
WkyCpCEHAvJ7zlb/30KG4gboSqCtD6U09LQiNDw30R3DmhmIdZr2DknZEHjh7Kfx
nDZ2B+y7pbywLiGLBxLMNCCiNKajI6PCC0shSMn91CinKlk3p9LiLkb67FM291m/
Lx+0rE+M97gQSy8fbcubdow10UyH8cAmBiXiK93tWqJjE5jNkHMg2VD9pkOsQvKw
Sqhmg+LxLHf6r9gycrP7qWSFEN9guer7CVzJbXfOdseDlBrT8VBLjYt+PV5duCCE
EHy2Zkh8gnn2DIqLM2r2epD0t7PsOjMCoe8Uu/yb1jYGo7dm11tpfbz0kGGOSHvX
ecTZhlfPQAWXpEM4hHmHrJhqZmW/+V9oJN+2faHFNNWpoHlKkPSOmx/+5U08mxq9
pB1ilnqL+WRM2M+2aUet/1WK+8kMbZcCtXDAmDNs1hw/m/ohR0NLy7EmUXuTFqW0
qLFl3KEDWHXAlufh9V2FmaW1rBs0XMzyO7eet3XfzCG7tE1pFB9yVQdzxEfEXja3
tKTMhtgPFKmvAh3VPkQQphU8ulK1yeR9HXkOBjchfH+gp2S8IQU+gIpk8Si/zB26
AH6XZWORjp7eTj97z+UhnY7TUiDsxxL6XanpSECTW+7jtiXaA77K3JORzo4p85Mz
ERtib5Zyl2N90sCAuZbZos5/mKYn/cxtdOtTqBvzXjske/M9orbzm6QVVvMq7SYi
XRrqkJGkQLTxKO4wS3hKIFq62goDKf5FCRO7IGqTMR58PsbuHQMgqORVEa4WMyzE
mtAIjKyV5Z3duxvxuz9UgiY0naClaTNq0CJ8X0GJxyUnhnT34cWwbFOvb8BQNrrM
3MFC42aevVrhas+SxFi4A0TPkAx8AvDLaftmZ72MdFru7U2EvHPJyMVFwYlPH1+F
UoP8dX8vsGQE9lUCtAXGZLFKrVexUqrHIiQerTYDYHMWlO8JG8QbTttET3+lNhCU
VRlunHLIBYxxMZu9IGLbyoo2K1P8dFPHLCWn8mvHBCndIZQdVcwqfCmhox7cU6r2
kl/pfGtEDIHN/7Jbzol/zBQ/HVUOcJ+6Mmg8MveLy0/0wHkh03KwoEIYpj136zdI
Yd8z9N3Sna6ocqe5X7Aij2h/bVPVv7FbIHjTeM0Pv/apXR51czdN5KroR4oKs2Wi
rGXegggzTkGi4Imq7sIpHe50szKLuAmWgq5K5ezjhwjB6EmGEGdxGdw6fjg8ndgD
ZxA0rU/JL7ud1BgDDHCAj2ASXCx/K+p5pyojuL9g7O+YZMvevNIwA1l43k+ZtMLQ
W8s3vJtUDGY+n8iq1+1SeTll4zn9kos9vMQNl6NfQKKfOy2m0Rzhw+UZB2HGqdE7
SlC9thJEBOj1+fFHQVvRw8eBtW0ljWV6UwwP3ZuMJ9BJNkQdpCEu+cZkRsjfwVrh
dcXrTMgyYBSAQT2uXikSxrTkLojIhglIo2lESkFc0ARMbEsMOTjFm1wRtg3UOSpx
74ooXwPUrdM7YSWJ0NRNL8pyzoqRyQATevOEcIVq01lA0mi7udyCUVKeNm3Bz6tq
ysi+7auODYDW/C7OIKecNeF84nU7zpRMcEenS3EPP6zleQ5BqbuKaf8V6WrfJyhE
k5dt8wdu+xbmNdeuTVIY1wnOzEj9bIGWSZeh9PUsy7DRGA4LZrYAgEcPrchh8uWy
cj/D0UpjMQGkKCBNhTi5dYgMtHZF8bAWdC4NF5cIaX6QRHcE5sr9pAfeZS+bBzxS
CwKNbb1arxpFeLaYkKnWLMldwEIh9v3ZFZ62Rey9R7GxnSyhwGuLE27ujc7uB9vJ
FfjJcex3AIO2CD3ogEK0k1US9hHgqRjytZJ5k4UVGvcdk9GJMJYyzULMZ4N5Wvyu
fB05Q6OfWGN75X49Py2B1TcmiyvnG8T6zthEx5kcqw0wejXCdX3VSiSe1yx7F3ro
M91q/SUEUVXKaLiIrxU3keQxTztrbmLlFAYKSoPfvl4zFKGmT9vdK8Bya/6yT3Ji
zrUw1AZOL9n7rvv79uLnRSSqtKPP0ryPgqGdywCCBE3TC+YB4/ZeE1HBbdwm950N
cg9ni7+a7EO1v2uptUrJapi9VSbDOoNhIhdeoybf5fjUB67BOLd1JYYgEHAOH3MP
QQJ9yovDNEt9uEvEstM1LNh+J8SD/0iyc+yS6fKvbMtysWrcZ2aE0pEAG7nOCMGp
cnnw2Hlr4+NP4pwW034RrxyJwP7xjzh7JWuNRZGuZglCVpNUn9lB48CB54IbDDB+
OiAyuz56f2sQ3aVhY/kZzjihECaQVUdApB5v7BVJeQKo+Yq6dnOQM3fF8zNPKxNg
AXaZqeyBKT9RlAWM9U/RhMXt2wm5MXKBf2hg5i1ZrCeSCe7/Nw9vdUZOwjGNxBlR
6D54ftAj3jRI3Fbz0EwSYWP7h2v0fZZVRMkWdctznlvZkdBuQE5kNbnTP0wDErOn
4E+Rh/ljO2eFkTCsd+FwqHD2RS6bCn+HjwgsdWITDU5kx0yVrD6Z6l8B8yySxWK3
z+bYDxNS2ipUigvc7U0TbldTDJJFU0lnH8lfQev9EUhywQ9Jgp7XPRHRtYylul8P
jkMcamzzOjojQE6bNyNH5HmwHgXosIXkJIE3PXi5GyS9RFOGIrdJO/JC3//I6Bz1
I2bkFKiV5VfLoyGIVl9Ebeko5TT50WH6KighVEO9oNDa9c8lv71YcvjAJYIUyvLU
sBx5MKPmNbn6BpxYA0B9EGCSdXLUwRvN3eZIizWag7pJ7peV6eK7AZmPP6H4dqB1
mFtqcV/7kpZbVlcl71CbD6zpkAPRJ9MH3GczzjMGpHVVvKz3nzFjV+WAl4NcRNbO
rCMMbTB//FPZ+X289UojOQZOF2368LBywf9uHvaMhE8C84WKBexF560xvSGWYzhu
EAG6S12bT+nuCmElimYhAqsv1nD0mwOVDdrN53qgSWnW3g8Zc6YcD6fZNxXG+mlp
CwhjrosaqiZ4NDkPoQa3+hZ2gTj+XBxahCgsydMxO+M0StnktCSn5k66s14119m7
/JFOjaGDLFqV0OMXhVizJ1wlLXuuYNFPlLhBg8RoPTegCOQt6TEYFpD3vJNQDjvv
/QLHzxTWWUu0huEgIZ03Oxc0K8MbsH5vLveR21roqXzxLAsfSoOaEyuu3ny1uCnx
mfXVf0yiVS4fvgpKZ/x7G9Z5VnnQsUzlGiSWgiYnxfOmGNlxwhoDRRtVUxiQxVqg
F4lNNaDf1Oh/H+GtpieiO81awpVKB5ma1aU5RpAfw7gUaAfYMoQQBXqsDQC3no4G
8BFALIC6hn8slBFsidRHxgv0dCszWXnvXCjP+MmCWs4v9VyvfZI9TffMHFwfz077
poLRBaXGGjUTGUyQUA9xeLDFmu8bLbdHDMSlEk3O7Ghpe1ueo4ZjHqHFVVc3rrmO
ZvVOYsem/4eFypjcVr0oWhwFXmwqnJObau3i8BFgltSlBpLUsORZCK2lGiHJ8xmk
6zQwCLdXrc/2fbMenLlwheZPh7UAoJ4zdZ9mjjzlTw+a9g5zsppYL7a5UKCrK37q
vgrg5TCNf3v+vbwqYwSr/LqFeK/GJ2B2O9qVO0pbbDZg6WxAlvtI5W4ikc2RPsjp
JVUNO49E83mMsrWfObwzHJz7X650jnVzMZGVuJHbqEBcbn39J1RaUoQqZ20Rr+fl
Cewmbae5GmAS00eqv3SosB+lsLIIfj6EKzFzaJsTIoBENDm+WHzeIR3zsOu8UpZu
DpbUnGezH/UnBx9RavpLq+mWrdqH2qv6mI5Wh/Fllsu4fJCBskvwZHmZ29tWtX23
/GpnSYac6BCMtbQyuVYF2XMWlEGNAzT6PUL6aWvn3jPlEd/gk6ncf0A6NrqK/70g
LwHRbALqA2j3K6i8G1jFUoLztzBzOgarDMoHOQKuHmki0MZTnxxT6iW77J97RlVW
j/ccxEfXuIovopEmTgkRWwTBYxVa2rlh4ZS97meOP9f3+t+2QJdceExkqrVgsam4
13uD6QuH13ucBze4CN2M8x2D09joimJnZ0vx0Te5TM5Z/7/+7zGP7bZWkcYUWDZY
Rm9nVR/Nko7BGEavq6VxCrd/l1YdslpkyotfDjU7fnRizMssPRTByrAypGpq5azg
anHunYv++h1EK+u7Fxa3aikGN9ngVbeMQWB32nCoZtE6cOB6mIAfUezDcMtxbE7w
79JTtBqlWs72c1QgjY9r1/V0NutWCP4alFwQLTf/rX9CXQXf6Fn521ojBYLY9GrN
iGhI8Zw1K5bAgMCJJJgiGS9Ku1sOKN/NGp78TeER0ELhHeWQ/sgGIZOFcCKxx4j/
Oq0oDQ1UBg+I1PCGvpJEckmCaylT+wfu2cQcvheNMLPRYWZCLuXi3RTx7hwMbCNV
4KaRAz5p1Z0wUGcV6ns68BO6eIiqOY+QP9tO/YAQoiJHQWvBL/mREVUSzkBSQRiG
z9D71eNyJnGJhJzA42Sb6yKyNljG0+hHhOYVthC6EhDCM9ALxklx7l7pNgeX8JE0
6ZKMZJOjX8yo+2UQaFkhpQptOXowoDIyvosSozF8/217Dc0kzt1kVI5LMGgrcfWW
nwcAMkGWsKAuVgGyOhMIdo8huwsOpNtdrGrCN2F+OqpR5KTPxD3vvvXMSR9CqReb
7+LGUW5Mz2c0BHZrSQcaUGHgYVEzCHa2kLFZ93KqV9Ct5udbfWr8kCNiSknq6euc
tP0bBWc1Ml26Al4/1huYxPCl5T2jU83n7PIGpBFZOLXMeiuB1hwB8m03PcDGml0Z
vMUd+xV2b9pz9N6MaZWNvYGq7DINbhNRDu9SC1/M5dbXAbXkzZgxsCcS6Ps3SsuE
/AQFCc8RWTBHiW8c7ioXDZKaSDWSfZoDQEC8yd5ducUleBUCUAcs4QNXkQpZthFn
uUyldQ4XzRJnaoK0qfM7jJaSuSrGqVgy2Ylqi84IFB1QJ6S1+lHHeZqDi6cOQP+l
g5qULgIPrwk7jx8fwJBmOHfWvfejb0m3v+5DXM7k8H+hwy5d2ib+TS8bc0/nAPKV
jkZLKpX0++8y5EgXWi/Jg0YdAWYzXmwhP0Wj+YEhO8xJhKQKrDybrl+AWpEBlGa+
f6BZLQTjjye42n/zgQTx278ZlyaTnXzS6GcsHnncdgoefp2wqo+Pc25xVRJvOpTY
g7xVsBxt/fD0/K9lAECD36xQ2tpiwknb+ym5qreP8LrYCTiX/DMZLluI5HG8uU7G
/8xtjRKORJFmvdYKFzR8K86e2icS39qBFZGgRzM94uB06RgJUGYvAfof5nr9lWaU
TL6UTqNncc7sziQiejVYOjAZQMcJKeYQKKtShxYF+HVcGamAu8Sn/JlBY+seJgiv
SWhrS/IZMS25I1WRgKyyzQT8ngqm523CIA21qc0eMlmA3b40BBpjIgRGPxewR0G+
ECpkE+8Lg1KvZp47LoQtu+usgj+GTw7rprhoCN3sXoVAMPDElizq/Cns5rSCQJg/
q5ccWegJ1w47Ri0rovqg9pWN//XsHCplT/W7uUd5bFmtaLAdf1Ka8U3zZmPTtNwo
J7yi3bGXhngGFjlYjf4gbohCeAACmIGW8I4W84DpAlEgUk1A/b29eouUDU69HL6W
g2+1Vm97OZXz5uLPcTN4Y4t/EJDcsAsKd2Z0nBsu02vWcJterlsDpJxkIta+oGee
a5pCjG6erz3+f6ErjOpj9TcPy5IPYDOsaUlkdb6ZNc2JX4hynY2JERVZhsKdM+kf
Lxau+AtSkyuTdQ3nO+4Kyi2gLnYkejANEcD0zvf3JsG4JQ87rHTCLiJtSovkrhKC
v/3vokEs/085Ju0T5zw5Ppng1Z9Z6RsQ2VrU71ZKltOvLMAmCwQ4dStXUyZxT4kJ
QKxv3gH2a7wQkYONQUu/B8rSqkZE9iKPDtJmO/nqfMLs2Ayq9mXxzPSZiIofcZY1
LK+RhyumQvipBFuFUQDOm/EVdd+9FOVvOhknrUJzKQZobHuW2QtvdlkgKGa59MHu
/SG1BX+Ioud7rkJXiiQHUoZYmKD+VpcY4VvSAb+KT08RMQyl69Dk6QflPm2U7VjN
gx0tUQMK1UIPiPb5FlRDXMQ6QzI74qyE2JPkZUnKngvYOLM92jJUd5yHRo8QBxma
VoeFlXUNsRTy9jsKc8z9+TewW2ZXZqiXx1brLXLvHW65Wk5D6c1gJK0kxO8kQlOQ
Qc+/SllZxM8cZD5TjbYLIR+5Af7bIM2v0W4KXRsiUoyB8POk8iU4rgOsOuTAvaki
oH9Dae3Nld5cHZRswwlnmGb56UQ88Me+IKoBX3J5P+blh19ELPrzI/FP6Hg/50uI
h7llP9Bgnoc2mrsckW0E6No9vWAS9KNE3Pi5zMunf1oxKmGOnU2aVAGwDIjgx6NA
0eY178hyc/LBo+1wsxxlbpVbtkRi5MKo1MAFZIpaVSasCbQ7gqCZ08kZ+3gvJLA5
gFIzhfUv4vpZ1VOm9LLv+UTAhVa5SLBw6+MYo70JFJxl+nH2X1SN1TjlU6SkhZqC
yy1/zqLCqnNKYq3vdZYLw/Eq+xcgGR2mCLjUvPcydDnq1DceK9rQVkt+CWh24cRS
LAuMjUe0QIz2WNEghBW72tZnrwIM+JqukijDEk1vg+erxZP6oWzh/uPo9mCTgxwr
7DvdcRBhVAHr5Z4iFvr8rzou7dChGFNKE3FRKaISu5OSH7OJbcUr7rGgfzR8ET6k
GKJDr6XCy43B1gRl3mZP9LOZDgYMZ5mzb3fZcooB07eCHSvItkhGMHGZ6oAKX7uw
P9XDqGNxQjnjij1oM0+DEYAnQRl1bNM3iSNjsGn1R/lvMhnnKu+7ZU2gulWAvyr6
rOXteJ0Xi9mZL3Gd0xPofIzleKNq529/FHGJuqrBt6VWHo7+c4jcOCcCe12ipZfw
iXLm8yHt6lOrxCjsN6MHosCuPoIX3oe3DofZ9+ysOd5USf0jyzFOiJpFRrW4Ern3
qbtEx0B3bgsb1gQdI4CaMn9xK3G0pWl2c1E05NsJNFCJxHzQkwYAxKlCzQiNnmzW
4InK5wyzJ+uSxKo5ePlsXBVRJ9f46w+8w8C5wWusyj7+BwOt/OhEZpB6AnpUZFnz
jwo4svxVUPyq5uNyH8wVxs48Nfwmmq+hm+OEREPPDm0wRwTZ/YwblO0OQ/HWeS4+
GQW8ri/NbfgrDDahIfPETl0KrrwqwGYoPCyc+PczYRC7CFolc3fx+tUHl3KvTF1I
G1+mlq+7WJN+WqnxOxyotVFJtrzyVGR+7fq5SJswAv+kXqnWmlVnmKSvRJ4RmAht
suqR+EcORkxei1DGHCyxBSSBg42MVaNyXJ2CtnmVh7WvkJ2u4ckerQw+YGZHL904
eb3Mdm6I16jDl4M02EI2XmNBYTwB91Jn++zfyHo+K191c6nwAlQ2K8EyfmbN0KUH
WVLAFQ6LPd1JCvgcyMiaM+6UtWVR04T4SbN/FI0o/dsQvm4W72TEnP7f7jIMX9aA
e0e73vKXazZnZP0+8ydNThlsv2EaaMSeab/NXwe7ZVbxKpF1wrHp/BQUhDLpkTho
Y0bFSviXvyIigAn5EerD1Wi0vAuIlEjYq5QJX3pgwkqE8rRLTRLSpUpt5DE+pnuQ
iaKsRtIXk9PIPH/pdU00MFPh+wgWN6B1X39bN02b4K54x6Xw+LDIrTIi+sGH6Orh
tgjWipfoMnPAatNihGkSyDWQZGfYr6IqycEHdC2NXPEwKhiqB/TB6yGH9FvA0tMY
q8CCaKtSnoXUW/HaT078W33jDjGuxdtqWVKLs35+HwtYqRZ7OjNyDY57JMmaau+C
pLhu0/Qu+zcjRXMp9GlOO4itY9/eNNQhLSJdVjoo72k2mmsi/KfLrVtWyrHmlU5+
KkW48dMGFi+jtjcTpL5/CxW16UaCiQpBKyp7TjlKwLf6DuyAHFRnVcKXw78YPzwI
eit+Pt7PRIkJqoTnaFdaRBjXo45LsiYOmCECbH/NMxaxr7pN92Vp5a3GcFLoAbtW
JdJ60M2f8jPy7FHp/2bIVvI0fXCUPMKKsc0aLBy4A+MGbTCFjocI1siey65lISQz
eEPiknh2ShSiIOQSyg3lnXh9zfhffaY3m45Hfc4jnjqLzUpZI39gPd+LrzOKxndy
LI+R5gRYkg/Wbzd1v0Bk4qp7cWpbH3cdvcrPWKdjvSCyYND1HLOBNpjTskPtXfhp
i83RLBqibeydrKpb3Frk+BREydmvlqDotWol2ooHcxi38u7LuEgVyRW4XuCCKEuL
ohwzdn1dIsn5BiCQiZs+MY3f41aTpUdi6iHJkR1OMMdTXTvq12giE6VdrtJdc3Wv
+NmTXVYayQf4LBHbsa4TqbkIKPSx5qJoz6kyZRU/0vd4OtjSA5g46rJde0KSXddw
hCmfHglVlcKVEJtoRwq0gnjfmH3CHpJOlMHLEsh471TYpBpyuozXm6IjcW4tiGQN
siT0wUa3fAEa9JPEeocz7VIH2HN5nIAZTyidkWYPtE6DptArxyj7x+GKERqpV8lS
HUf2MIa6fDY2zWhZCy0yeXOyQOYAlXzueQ33PON5DgrUfrie/jhz0hiiQdChoI7V
kUkALWH/tQqs/ty8etSwMF0aFCTWDWgU9avPa21EWlQ/MhfTUctcBa8s83lO+jQw
qCaNdgg7atB57UWDUq1r4Xc/e2kjk4YQLsM+zS6KLXzzSLa/gmFm13A0+WsUB2Yx
uqgKqI5v86gjBrz8rGROJtSH9+h/6fqRY45UbBXNqg8xKsbGHMdIm+w92d+1+0t+
0AcVrJ2ei29pIADiqWPjottmXwMoGGUsKWdfQtDoqm03PB2sAemnd4qAW3y5cApR
jfKW6QFPPTo/lNlAbFG2AkeyTwg5MPnLyTYbNDcRsG1n69sGNzYfVdlT9bTOGyT5
53qCNWpeDrNPXB/+WJry8opMygWuBGdSdsvlHOIBi1OnGExACPMROowaHibUSo4Y
0om8Rgx57znJzjHfhKKU7m1R/6AoBSa+iAHo/kh+mb8DSQAt6dRL5R94UgZUt17U
Iv/vf/mGc8vk51QIxUvni9EpuRvwgNDnrUOG9mLmDtRpqfYmxLBzq6/qaixffVN4
eTKZX3O8olIEAEcK2OuJ2nlyZMksz8F17Tv3U9R5t0BSDcmoasa/H0agEF6ZrWec
VyVRkF9Eb07JPlI58pHpxcn71rHGwyVTb2SFk7aEXcdomTsw00rikkmWLEogKnDj
FPJB/0HnuSOVU3XAw2DD4QXLXJYW/QrNHsTrqnrAFHIfeskWKZlHL2w2tMGinfoQ
wBhYJPCb+iS+JxMaU/I5qlpMoqg5aZnNweV1uwJv4SlYi+iedpImfcWokYZf9TSL
qZFnxuriKoTba+VzgSPEA+S7PHW9eN/j/6FZfe/zjDQyJehg/OWtiSPP0dr2QMcE
icbtzHsBdRBXEXsGgb3Xeu0VrQe3R9tlAS2ZtRCCf01k17fRk9343+RBv6JWBAGj
hUqBbCV1L+gDkCWh2yqQ/zpJCn9CfrLygbtonMx1OoD78XN93Q45M6LdB58+q9Z7
kFoVN9RCUsQFzX3ly4GC/RZNGiHhp5rye10TNAOzm2pvHFXLCus98N+aN6MgqKLF
5fQe2mRySxXB3c1aIYIxEfQqzo5cWC9xiXbTDaYxnkCM7CuXIK0XWjX8o/szA7O8
ZKZ1fmLC6yQezDiUtrnjpU43Nwl4Y50zUBmVSP0xz8l13bel76+KcGpl0QPQAwcK
LcE4jYNKE7Gse53qaIAZbG9n9+rYmfKfZXnW68Y/cJSBskEJH0OLCZydM8nPWfkQ
WrrJixrW4wmK4d8pflzxOd2N9T4/lwC9iyUhs94Cf+2y14fKJM+CaUjv+7nAWTrt
Z8uF6NMUW5E8jeGuCIrC/VVpgWLxKk+7QBnfvEECGjsF1Dcm/r3aFGeOx5HEIcbY
mI/uR1KRqYaNewJByafD0ZTdMfvOV4+6kVL2H4K/EnGHIt59v1Jiiux7+UC+RV1D
2miMYvOyMz//ofDe768v5QQEXZRXMPZwa31p1/mHeZrf+kJIzDalc0o9Q9dhACfM
JsdBPb0ukBPHBUJFNQ4tF9KcRiD9x8dUxvETzyQ66HIkcZaIVM75LKZtDeJXTrvi
5CzzZ6wHc/aYQGTFUhBHNpjUY3N4YM76vx1QSI3/FofQH1dmkfInrzxJjep1wLFY
rFF7g0Z5Nhtg9H60+Dmied8kemJ4B3Pj+cPugLdW6xKMYY6iovqVZ5J/u2k/3hJV
IeDbmEBHWCkgSVNHp2AG6eps7Wk8cSYVzEgHGOdzrS/yCxJ1JVsyYLMaeyORNIRV
75ZR/rwaqhEZPuskZLCNphmEn+S6ZYJNsjgAOeONlH8VwepapZ3pWzBcyR2+RyOj
VFXmjTP+uZvhPWlcepVfQHDlike/ArSKTAQYZCQqaJyNnxSenYX/a27/q1Nsz6Ly
TVTG+7YSimEs7Lj8GCLa73QS4uYXm2qEtMdFNw5OhVb1TMAbSA1Q3MBkAbj4rULs
9CKiMZJxURGFZUU6cJphnfnhfk229dkofoi8hyMsLeLBHol6PkeieKab6Wyhjsny
i/BOR/umMgVBpS9Y4XiO1i+XthYY8j0WhUiZAql3t1A3rnvSH2lkSb/Ow+lAQhtp
1Jzg+6Jd5BjcUOVDT2OE4kbPxDkQ3Yq4YAk5Bd6SYTXk/2oz/vSjFGYZUBto03ZQ
xjzs3EeO+WOcX8v0j5uIO0d9G8R5jTH/DvQvwq/Ge6lppu+etc3vW2CbSL8dlQ98
3jBFz8DCezE5Pi5WB1uqZzwWxNUsm3eoyQfjLHmhmY6rcBHnRGX++oTyL0z7kYKZ
S+afjn6T7f0G/BxvX2pyPhHqWUg1m6uR9Ro2s7uXS+Kim+8cfgyXzE3d0EuGxV7n
+VTb5Ab/vuAuiNvrgLQ66D1zo4bkml39vHERHrR+f4Wj2XPRBuDnb4+XRynDQoKS
/lzwW71aJ7UJKqdKT++gENlaiEOHtYmjndLirM6pBKEepshG+x4PiquqIQOTdjwv
w3AMCHy1qz4B8e1VgbES/YCoq+/Wfat7q4rQdDH5gPs82XSb+YjFa1SrZOCROrtS
5Cn8KDWAYEXBaJ0ZDv9O3ax+Gvvj6WBzc8vlEUnVqvujK/E0vZ/VNvzgANlq7xKk
VF0RvPYfj2bE9D5/GmkCpke0DjhNEWMcO1OfjVClVHPLqxdf7Ecq06jGi1V6njTK
CeKcuyzY8Dn/jcYk6YKmb0/O2zr28XwnIaQ5/3VcQRPpqr6f610GpZwLigumyB27
lij860OcsCXO38xSuivaJ+U6cWeXGVqr6oITixrBUR2knetTqAM52Ab8Ld4inBAh
4V/n5A/0NnBdO8n5JGdIGqt0FhC9w6bHMihPz/xwPR4E5AGEPrOI2Pixv6O6I+P5
uM7Akw7rf526//ms1Pz4oE45KO3xH5G2S3w/eLpJLBMRv3X5HKqn+katvPPJH3G6
4scsONJ0SHKVMA5lJl3otSKVXbMDdXtL0vduHBlEMfmj8il5yEM93MRIqDuoa8mN
kT/FQaHr+jK73uOngfwtDWz/CEDhADIBOsps5gO9kfPziEo1wIANR7WxZC+8ARJ7
ertQlfTeaWG/8YbFf7Oj4qYZwLWZNSa+TYHLhsjVDvHpSh2tAgh6YRzRB/WEe4k2
zKbLyJAvEICdxj3pRXMTI6aqlZBFKcPz6d5SD5Ws/LxMQomO2J4PG/TTBrDu/lEI
S1r+FyQ8nEsjYdasdETdy57rCO5bJQ7AeRMfIB4Kj5UKT/Aa/FWon7zWFxiZ/d6p
+w4xW8M9nCIaRUKjUizJFwPVnIz1yp4VRRdzrIvUYt6BZsfvOjTD6SsXyhUALvg6
7iH1bH7qZfUcBQSL5WlrWXlLFSaJJ5rxgvHztSC9dmIwJUykCpnd9alLB3BNW5ee
2HAs8OzGLggsjkNj84IZ3ZbC9SaWPuG53ojKeVCK//40KD+hhGesWgnD9p2qRHJ+
ycr7UAi9Ray4DvEO2gdKL6fjrPGKGfFZs9RvfLXPhnWIbOdNv8/KHm5FsWQYQVkV
tCvujWNkUE8IKqy9SBG7AmZYyXcXvcUCjVleMjs7qCInrOTnO3CdakdV6ABCPaRW
9QxRRPf8vxcFWwJeAuQROF5eSIe24PIYqfNDCcjktejpAQuYKriwS6xER1Tm14gB
V5d7MHUSHnmqilvSUtgEu20obZUVqFaCtWDiEtM/hlTPQlyJhluZKAvFW9+ojLpg
fny3p9HyHX4oYA7IqkxoM58YJldbTMbbd2dnOsEefFdvk7VkcMZvQS0LvUSGMYnr
H7m/LAhiRGyBxVV+J/lACaAIUekpvO8EuuzjfWnklZLdgpxKc35Nl+DL3FJ0+eCi
IqF6T33VXv4Z/eg2P3O/WWwY9m4nNkPEPT7Dv2Ece7H6xlRMU7xEA1cAx1EW0Qkx
UKjpeoacaEw2/vEgDMVH5f5JCNeNMyPTOPQ3v7PDbe3wDYx19FGA4dQnB4dgPhSA
OIB/47xiOOlYd+xcRwKnaatxH/kJOlhTBridhlMNNggkyOSctKhfSN3Skpr4anQ8
fd9SqaR1Skrrh6o9IzYjx1qYVM5pk+5uoDUVyFHcbn8CtLRQypne4bETfQulFpQn
DVTHgniX5i9lfHeh+x60st+H5t9YxwngdUeVIjX1DXcWwHVWelghPPezqxe2nQxt
72zI3iBlWyUtG1WtZHx1k+lCU0tnRgofrBskRMtuj8GpYxxaMmQOp9t4ZWXpDei6
c+yKiNi0N40QpYxMQ5jsbDquj+ycTOufYeMrAQva97f8KwyZ7zTLZUCBACH3euUd
Xp9saU6lhAwxCZ0Fwp6Tqggak1L9P2lE/zlXNolBFn+UHrtd34FrwH3h3YQQRIM1
bbBVZgI9J0mDD5jHKCQQZjxcpxeuRFlBIY9vKkd2LlMcqwn0y2N/u+f9OJHh3LYa
5le1TzXvI3WgW+sJ9xCpPfKB8772JoBL4QM4bN9y+TMY6gqrwDoePdFIufbm7gA5
zNCavApEeBuzcRQiI61iGmvAT3ZQf2sKcSdqeWsLB75QuJBHYu2VqFapwanJOq7B
7HNbdpfDhyKX0frytp/wR1H0tJ0F4JDmF0UinuiFDSusSzRVEfNJ91EVdBGFVrFe
Bq+dLf244TMvuI0IYGW0LDOOhHwL5JDB8jjqqj5lF87yjl1wpSYyq8DTb/lhjAal
ThSRVtFHem7znAaUmOl8E/B0q98Qsemjt0C2b9dxhRsRF4SJbd7VaMzdcQuBX6OT
qFMCmgTQngAAJUXpuZ8Cmw1C2PICPCgws9Pq45Ww/9Il6RQpxtFPNGAyYJ7eVHuv
6TiMKhhE29XCFgVD938KcgwayoUvwqrz9zoR8xANqjjtY1FK9L+QL1MFFo1EQTC3
qawxoIlv3gAK+stp3KpvBvhqrx13cEzuu8ZBRvacULRT3p8od1KOzOJHZQbqgdj4
5lmr38LU3XiwY9LA3Q0JtejI7TPFI5b/4rppyjuuxBsb12fmzbp7d1XQByrQsWpu
bsVCYuW9mqru6/0d09l0q4e3g8XjEmVLvs8/Ax0hBuHxbeJvIPr8loJuktY3AW4r
IegtZocG88fd5ir6C7UVNM9/MFFFbuZxRW9pvN/b866Wn2wFuGgBGpQHnT2184Wi
ElyA+qvIroJbaIQASX0m7uMpYAbQqYWxu/VnyVTyeVvyvjOW1fm8q7OSvm+RYInQ
ipl7beKY7d3U4zIiAb12aucHuGnAIpPP2RFqP1w1OmtGnHuZVSEd3vYiMaEB3Vcp
+Lcn1DKt7Ut5kumMuiPOvO9fzb3VnTJ9+9Id84sZzlQ848DI9i0/buAYv1QHUNUy
35c/TBlblnAUgISv+ujazYmPkJvE9kDhswd+c2dAgbHxr17n4LSisGoSigPzgZ8L
xJtrzxXKA/aKDeXrb45Rgfw2BcnvUNodmWDwPT2sz/fwINRcRskRk/0Q27FQXr3u
jD3K+YSwjHOL+w6QktsEgx/Xx93GssJr1bbghas8IM5yzJ9cilqqw6buvmC7Qc90
d/yk0VnNF7Di6XZ5e/MY6+49B6zJ7mEe7M8cyArGuk0kYxHXrP5GLDdldeu+mz1H
uBUVInStklcNpu3mUcg0jgYLzAG5aqZdRH3bh7Wtrp6UUKpttR2IUn1W2HNk/Fch
prdsVz3YS5Onjo1C/qxFRhORsddIE+CPXPLR0B70aeVQ13xCvpqpL5LVtpjSqwoP
P2c/OHHy6GvCp7zvYgiBycbxneVLKLqLX/Rn0JxWJ1viRVTIv+BujWt6HwsPAOp0
s0ikx2TFujtRewu1c0y/3QpM/2Ff5Qx0OvnqLTrMCUgTEi2V0ApJSRbOe1w0sOC2
y3VQvlpNrthdFMIGJRgdYGV3m01P9BbLAeh82Alm1XDGcRyaXLB2nVdhS1uSKZud
Q/xrE1OUuKuvQdWvCqe9Y9XRhfQETBL7bFfxZAupuLYcaY6NTwlGVpD8GTmUaeib
7+9Guz/OvDk8r/zlJB9hbdvSGux9XTS+eKr5mQTgkg2Ddh6dRyYhduZFnyb7p0mJ
tEKFxzVopcGYQI6R6mDle3UshJ4vmwE8oG79i1qxah0GbmYeEbT13VMi0eZ42yy+
QiA6paPKFVzItoUOkIpZfBpSzSkW3fH7U5wabQcJr+psk0psFVJu02d/UUzE5vOK
EVp28gpYZMFdA1hxZYLLSZPXk/XZFlIYgZcKAxSxIJhY9dRCpXFRbFoAqNsBrC9g
pVgcJF72IFXvbM9IFvd3R3T+NTB7yF3/fn57eDFMPyc/p7MOYMjFmTpcDtR4kYMJ
jcsXAM68+WNI7oIZ4rtNiHOH2D1OlzIM/+GfIgcqXMLf8m5n5vCb6ftF3Gup18um
HOT7LGOzC1t8y4ZiDbU8rlHw8+Su20nN/TcvE9GI/fXkC4HvyAw+hoIij1Fvz8+G
2Cy45hu0r1YTBV+DlDrkmb8DVlO5Boh9ZZMMAAB2sgKSfzqTDF9ysCK2hp/qBNLc
5/uUlmwochaJvaUfh6G/xVemVPEvLa1dGuiLGmzptrm+LveCEGfbS56Tt33d8Fl2
Bui2Jo+ySRJn8lcgxBdKVmiaeCQO3by2L34JONoqqYMSZgfl/pYbMkVs/4Za65uu
lnOqWooWxdPbU4iVcxZhfZS+7ez3Drq5Wz8r/lZ34mrW71sPlc9IxODtzUAHxGHy
TwXXQeoJURoZFwbiaK/sFfvSJ2Pi3nS5QZ5V8PmGAuMkZYfaHxg5FKcVHYikiCmh
W0SFvAzl/vhc9SHxv70ffX7LBuVk+8V58sqxi46keyE+Fsph5/VqhzsLj4TyPQnJ
ThckyvQJf1980AUeGEjNdZiDP/gEwJhQkJIqmASOhj8vKm1DCRIiiTmnUwn1Nmaf
TtFl1mM8lGrb8FryKKY6/TsCQl8MDwDNg0dLardy1DqkEKgmhQM4yNdion9Qv+QR
tOqCdApj7u5Kh0J3JraAs5B/CnWm5a6mn0ASNIc4mOzwlNaNYj2O5bX3XISn2/Ya
cUGN3RsBgN2XgANimbQ/4Zvyk1ZvFIdQJIv06PkKJdRBlamoxA8Pr1wa6GOjEkfW
idh1qn5HpF5k06d9ROrn64DHpYATiiC3nOGz4jJH9rNv0Q3LiW2K3msEydBK/HfL
R3fSv8X+aPM2pUOwpxPrT6YUF8TuHl/I9mjF0tBaB4GCQ4dULVMXQj8G3Y9YvYjb
pozONe3ghX0lW7CVtIZdGqHRWfyW7pZ7T6mOYvLH4nQnloF95ny5M5O47sXtY0Fa
j77IhOdMKt3SrXErX0/iZ6lqMzO53kT7mmmyKjKEMxxOPCrR9+8vDuAmk7qr6cPM
kiN7PLDEE7kzkQG1qhVAWlfdSFW9eUhDZusP+8LesQ3ykSGGS4NuUpzrqlV2msD/
dCb2f/iCq+6pY9tKPYo0ysHmtACqwpgsvmaUEM41HH2el3MA6Hn55R9j2IYfi/qm
GWDwjzk1mj7zvoNoC3eDcE2jeHq7ixjBZqOrz8blW7dQETK7RptuHciW/5bqX8/p
k3CUpzduSCdduPGiR1IJg9Rr9/6rhQ3rYp5vowxQSiRBRuLlRAqveNPwvDYceVS6
DWERJ1F5YGdDio8ePLqi8Hxq6cy2GYsHNFHkLoVLx4EK+qtfaNJAO3vNBp5+6U+6
r1tmJcGhXgEv1LNdpgQb84lRrZJUWTI83/gneDlYK6kEN631Z0v+Z8vhEYvusZP/
zIwyOswXolKTbf+CI3W69BeywamcD247uQ68RjIGcm5Xe9YQqKHSlZJM3ehblygQ
a2rUSBgryGceHhHzyzjv/S4kVKNFdE4/6QWBQNzBPGF52xgxVt/tssU0STTkAG0I
TjeqE74pod2eC0DP5UytIz+6ZYdQUMYrb5sdLx3cIDttX0EPOocIngKsXAyufyg+
jkQRmJyRL13xuq8fXxTfy8VNoLyLTa+/E0nsJyBwpqyLvkU9Drhr42LeL+p9SPHU
s2Q8jwfLBYCpOusa8Y9Z45t+8KDaZXap4XpXzUYSfdYzM2x/jFyx5Ll1DkFLn9yx
6vIIsvYFIFUFJued6k5Sz+MvSlq8lsDjUZXV90z8twQAg61PMRWjnqJKILIlO2Wy
lAqjbVlTv2bOcmUP2UTlnkX/d+xr+Fri08gxl6ddG8glTrzBV/gwf30c6mRFqVc+
TzvHM7Y1/v2jS49FdILUGd+TXngvPQDNiBoD1C3uOcukzlFl+Y9Tys87Q658tH6C
5O9RPCshvN11uteapjGK/u+JKqwO7tLOzbuz2sldHtkak3qO+SFxgoOSF02Dea1c
DPFhSw6CJimdu+/9DV3uR+Ln0xBGHtr6NdHT6OUxMiNFBC2F7DL6lPwMnyVy6S3W
oGIMIEvdye6cSWWrllAa1F+G9DPFurdk0WwgNffakDpM8WMWW+ZKy/1APqFg7cbC
qJoz97ivyRZ+yqdB4CEA4myZ5A8IyMNXU7Uvlul0+DkXS5FNhiuQTBHINoMoszBP
J8e5ZRhZq3eeClMy/Ix6K5XMpGJ1k/mCZScyYZaSnLgIR+9C+3k99goP0aUrMTuj
KvQpLehy34hPfHmeK0NVeM5e9Y2ueBQfxfaJL2QrOpCxMO5qfFBI/nyX0EmIPubD
ztP3mFrEEFIAG4tqEoNrs4X/xK3PqaVhDXO1RntvxFp99J89vpOfTRF68nRGu2po
ZrygN1pZzDUy8BMS7RPEFjae9i7B7FVtj4BHpkV81C/EslR6eBhdrq7jeezyHR+b
Ekhxi8HXFnWyMIEOdQNX36X1QeyuqrjoqTCQmomixJnIothIxZGlVoml313vc7l+
iG68y+hgwVexBRtCm2HlF/iUg2e1t3ULZAt1e/g5Z5COD4MpRK79jQqMlByvpb20
seY4rSFZQc/il8RIlaUNmmnPpYozL+oUFX2AjlUMutRpYe1gcjrvc8hHmea0qB2M
fbgySSlCI/7g17VTvNQ1wKZ8jS5TdGaIqU/c+Mc5zEn6N48RKZNmbQDI/7oXmCYk
I+gN1fNdfNSaaEq/LpNcp32woX5wHCz8OBz4azUmhukHCKoLhVHAQc8326JjloZH
nAZgEhsOH70nUQL8oJrcf/YLY9eEcVXmm9KuSiXqu73GHXBVEUtZdmRFLoBNO/wU
TkZo/8qv5aYhatBnVIeBtLweWLAw8RUnAe+cdWFwUkX7ckGq26yFxvvsJZUocEyG
+51M35qUrUrL/auhCMIZc2h55p4i8pFB9U+BHifNaG64HuoA3eugfJYSdiv46Ppf
yicMpNH3My3uBFFxu7MydRFcODr9RM7iqEiESrLXmmDBFy8oxXFMYFx7zeen+KES
efdKFuCXbYMyXsEDNWOQrhHuBCENIoSvjTvRvgDs4+NQdKe8x1U5w7AvEvxqe6M6
Jf/4WK0pSohCGCBE3RVCPxsy4bjg4ioElmdgz/guXs+Lwm/gWVHd84I2TNPwx9b8
49kIYBRxvoN4zS5l0SPjLnrT1mk/QqwDakiBN07NoDJckx42bNCJngQ9XZeFsUFq
jKdr9QsqJjVC9BKJ9njrC6I66AC5eDpOfLpaGdWJj+RZcky4gBNx1ZiJOrnlOs2A
NkN8NY8Ne56wyNrlsNVH4y9zYSb49D39/eHmXXtVHstq/1wLF4DByx4sC10j7W5t
M094u9c7sMgStF/YL5uVoofBq9LGtuG4PCHKrbDP/x/NZu+xgeuDNit5TUapq/SS
wNFOcBBRCEGmdGwfGvZPkd8lLDj0bnMVdZdxFAneqVWEVOF60iEEyJcaAPXISP8m
/7FTvU4bI6z02ivUmkkg27vNVVa3FJJUWqYzMrRbpUSX25lmva7UidnEdtxJwNLu
dXdTi0bJw8k00KZZ3NzNNZFCVHBZtvV2XXHMYgFUwMR/01/iYrKzNoIvQR85aUz0
qP++SRDefEzLWkOl2KDHgE3Ui3F3agqBW0FC8ijGkAAZS//UFgFCnkObbWm03+Rq
thvHbZZC34dfmRNTWt19XxOAQ/D0QONOzIEbpTGNGz69fxgMqywN+l1DSF2FSzRI
5AhAVzedSu+JbQJ2QVAInY4IbTglkj9gaIa6wlji/wIp5iYakZdWrpFcvCE3lW5l
SAI5UUy7/L/lLWfvTE8vTN/uVsnGJQyEtoq+0Ywt8m0xUzB4SmVuUMRb8MsCjpYp
z8jo+lcvYymV6nSiWpkaBlU06Y8TJMymqP32wWnW+YlEU2c7LXJSR8Hd7R+WJZSI
rSPA9zevHMX6V+uBJzldGntLlx+e583+sruwjZdjuXlvaR7HlkLgURSN5n4uWQB4
FSFI/XTJJ9dNN19EQ+xDSdSDErysP0z0Rovd147wTENwLMjOgtSUD+8m4jSTdiFQ
pn+5Hi8Xc4CUmCI5ersh9e8BK62U/SFktEXx99/PZk03LNIubJchJLCZB9ealK9i
d8VSvp1Ceh8toa8PbRA9Ux4uOvJ303MKHQWgRsQBetpazGD2zQFRlSiRJpqoDfMY
eZT0KFiDqnUkg/giqvRjqXYYAj6ineRP8+KNCxvUHjkdbAUJVftw9/zBEcNAXg6a
xYLA46klRBwcJCizlHu9YieWMoEMRJesnSO0vb0Qyt3IHKO4AFU/QRtScNeg/Crn
z4CEKJbYFoKXsNporkdukQpUBuZAgO8gI7Ip1qbQORwaTuDW8qqudZpuHx6exn7v
svZu2H036CYZA75uG38rJYC8sG8POwlNaykqCSIR3ERVxotsGhred1aRaW8fM7lC
YWTmTYqqP4/NWZ84kWB3gKoMkzAG9jNF7IWZKJFWQEuhKPbDte3ELxHzqX/QRQEH
0R/NbqUsOiFSJP3Sn6xTZoFJkqQKWoxosXNdUAZZvNc+FzhrFZdIdDZnZ+95+JHh
iwIV1AwDO0+UiHs1921XvBNq8pVQT9dgKvMCZ+7SNkDJgF5LMx4prstzgRiMcF77
H3bEbi2RZTcAfk/Vhe+0ycGx5hj4iFEsPSMNBG4Ul3qA1GoZm/olzE6Nmv8xY8xH
D8AfQ7+1dfKUZss70vjTBLHcnpOuC7KmA6JA8dOBXQcAkB1N+9hAV+oXE8YEeHyu
uqjUoF5fOnyuuRhI1nryZTFJKByQiOTNNV4R+J2Z2bgl6H9+KmzygKrPPQdLHsIk
uSbOiHBlhtuDVxMG1rj6qzKoljwDl9XkQbGFTE4U+5X4FrrFWFqEB4UMlGZ66sFn
c2HhtPjF17O2rvp6hieGWz0UHHoBmpaCygxFraVLSl8CCDvwdKc80pIkldzD0O89
aG05Qg9ABPYo6LJjy0GNdKf3ka8MbICgmS16iBB5fsppimd2wzX7YYnukiR4TQNX
qwJg7CpVXRyCyc16Yefkd6cCxES++/+rLVbDHUAGJqUtLKAPtBNfRRfuJrCp9uIi
skYuo78cTjFFDwi6qKrhpE8gWduk5Vue2OJqWk6o8vVKutsPKLZkhxD7AxDWmwKd
bBn0cYAp9PSx5ddTVIXu6K7lGmUbU8/aePpaoEbSTt4wzjVS6z3/ZZ20FY9gTzXi
KO9kIVWm8kUPz6hQNOf+KhtbstN+5aMEG+3KmafEgEGpC8YNdj2/VxmbXbZzTNpY
h2jaNJAu20qqBL+Z/dke1hpG8V+c7f+9+C7IUe8sx6ULrsnbTQkQkUxbJWKWRp4u
EBvuEFiEZsIMwHBtT9xsyKrpOlAGWWwJVD9t9HnmhJMJn2VS0xG92jjGAp+nPEF2
Q0w68n2HE3BvY5/y3mqXmCGKlOfO8H9XVw6nVvMhkX5JcjI06PPu/kCwrSe2vvFg
F0XTvwZUjvgFavvuaiE8TrpCXWxCrHXD6ObrMNHPx8U7VFBJpCHkbJEQGn5iMcax
PGLfJ6hKbrQNIPAmHTH51mmA2Cxww72CL0sM+GtneEEFOxl/dcCszt2kLkEnnpUT
7yUczYqqBIzEOzx0UsUdknYv3yLu/VBQaJi19qeMCarToXA9LUxY8ecd8NyGadkO
KgkMsVcRkNa4+NvhfpBCi1gNTHC/UZpIOH1L+FDjuPCoeR40ZpX1FQSumYyPktu6
dpsq/N5cesA2oDfEBJYeTpZIVdsC4iEmbWXmMpFiUB6PTdRPST/Bl7SUvpm5W/7e
Xdo4j/yBA+BmOSUmXnz/sLdPuAOXjgvEnfO7Gz00gfi5sgscF0yU1yJ00oTD68qn
FL4yMznq0stojLNGnHJEopbPxDZKfhWiVFYGfYeCohjiRBwZ341QVyceBIr2kiK0
zcqmsRuko8wRsZwgu8wUNny6DTqFPCPEQzbsPDZ5mryPsx3FFbQ/USU2pes/WKw/
JViCV8oP/8//vvR1lG3WNsNY+hQrLU6GwGAsEirbpiZZRZzOtTdegG17HTNepWcV
2pm5jf2LdBstO496AGJfYtHPmqhLFDHXNPylslqfDFyr1iVPxOB7SrgEcBnRDrU9
OVuON0wcEGFw869CWnp7XhFASRdCx3RyGf63RKJK2GDLxrr/YO8q2dRhplkbkHGi
4E6WcK3rc+E/4KcprO+bWLyiybCuVcL/luzLm8jpChr+owBw54/UahbHHJQJFa1+
P4nrkV2f80NDVRoftn01VdMrVInlBhy2uYk1ubBh5UNhZHNlrukrY9q9zUpTgz9r
v6qAHLNlZhndiK7+9OOyoOa+MXSEIADuA4ruCOXhdjQ8HNbBbbdvbpfgwHIJis8n
cTnMkYjM2bUtFYSPdS1biskx+QXrs8leK9ZycxLTOe1nTEWQz8mSZKpijc64dALE
ZImGLQlu0gCdY2h4B9fikwOR5dnxMXya4WwimaK6aBal//Nw/AmKjIizjUGVeBWu
z5pyeZ3eLGQ3XEgGtUIUeo0TqKQQBaxqIgthVKcGwC4SY52DS1eApQpAR2eUju/t
aRo2C1+KgDpzoyG8+1aKzC3yN/6/FcMeYcpCWGOn8VIAjEZZtCEFXoWvuGBS6vvC
RZupkx+vfmKuDrM2AgmiKhHwLrz9blQbCbu9rryXj8A02gsQDkwKgA/iqhPd+PrI
RhoMjIKajOsstxFoklsJldENcGVwfYUJmNT3/vWtNVpVc+YxF3AnKhiVtpx7zDKQ
IwHq+D/WorKa8EjxvSSKkDlzKhDRwq/UVqkbNG+00F3HfWCKuGgptgVFx+qq1Gel
BDYGCzzmlBh9hWkHgHa8RYUbz0jDzIIsYJct7NwIHDu/gGcTjrBZkVRlOVbXIBiG
exIyK+gpvEs9bucn/OqGXz+oJ2Nd4GxLORSiWuLtGZ70t80LRXQ+t3j/lHEdmtR9
n4eoPH4vugyLUlYvKCyBXUsWnvJWrAoL/7bdoM9vAEpbIrvJFsRf+3bopvkAWtHd
ga/VvJum1KuK7SH6/XiR241Kucc6y57x5mPJ2SVsI8e0FZH3Usc+t1Z3c9hxTTN2
rciJK2Lav9Zd1OCKPiphgOhg9Y/2EY2nbBANu44WlZz0FZBLm+I8V3e5UFfBj3ee
Sjj5QndLpvdRv/Xxt7mWwqIUPJW1reLv0ZxHpiM4PU6yOcSL3LRIsYvCH8dUwnEo
C7Xvu7Mx4L0xLgjIQ6A9hv60YJcrgpYx97JJzls9yKS1+7Woxg1kUbogxeR6xIyc
Q/yIGxCdZtjmGsrFAobqAu2dtKQThvCROfkwmReCaQ6WjrbAER61CL0NHi37WUl8
0pvScK5eWijVGiFOqE5EexZjVslrsiQI2CXaF4W7JV1neV2gGR1Xnk9xVkQokHZ2
o8X2TKUjTAZDo6r7cMZ/4CDhjieMnaDY9KN0UEU5zmfuAdDnGqiTWCFZ/ExA+TPz
9KkzJQHmJ5PX2k4B51A1awp4E4XD2zUnX4dnjRMdC0GY4Y4xf3I3NscKL6MwTS3L
bVKlbCZ3kijwlDT+zPrIZ3hhhPp6rjKxZOBNts+msr2cAgqo1rItGOpDClTFvKs6
udGBmIJk4WpmQfH6rXGmmnkdHJ4cuPcy0rx1gyNQUNFpla8u/6uGlo3LOMHuQHie
VSPkxD0gL566pcXLPDWlrAT5P6IB8jdlbhlKFd+XZjI7UOzqK12VnbEjuqgFxU5N
AEDeDsklTFJqTWTffrsMJrP3aZZVcy8ke0M8ah48KDb3TUOI8rhkRJL2oN7VJCVA
v2dEURxbg+W6BiTKfjKgUSA3fKBxpw+oZTyg7G7PAFzIFnvpPPphdBc68ihBLdL9
OURt7lpvD78wwj9MjsunMYFWpjHTHA2fAF3jynG1ioc7hc62r2yEHmulC8TGIK/2
tVLx0IXHDGfoIZE5c9Eg2Ua41DOhfjWxYYzUCnnisKue2EN02zOwGUdjy8P3hagO
PorOhNdxTUPKVwqYKTJZnmcdGppx+YP0woMhkeFAyh5XKRpRofWv4U/MsDhDj28w
/6jp2B/cCVm3No+NU0e1zSaTlwnrh3tZ6DPWp0OSW7IVsiocwG30coJvOQ+K3WuD
i9FIg1ur8U5qYk4qV884ebL7Bp8orOz6GMVqHwi6s6209ThlATifgADrPYLkW4Sd
t9HPapOdTrLqMv5q0nxfOgA0o737mysVFEk1pdEQR2vJO80dKnc/Cqqr/SQJf8f2
p2xIrs7k8aIn5Bi3x6LtjyvJU1zdG22H0nopHkKbHuqICiJ7vxD+Tz24h9U4NPy7
cm6GBHRLinHRu6Ft+0JcXqeTkt0yp1nMaSTOxHLOJDGF38coyovp2s1wJDDqF0GA
lfbGp2+mGypiX62sbz5hjKSwrxNUTDgFgjq+ARcfr07VbiYNbkIZVt4MZbJg78Ts
kJd9PCMU0tSY1fK4OrlnPF1OL8pQ+JjsS6E7LnI3VlBkL3MUaChTzb48aNvdoVwJ
jAMy3EmEhC7C3/pBMkg74Vjv/IarZX5CdavwgCPlV1+BuejaKD4aXp9cgMdxHpQ9
mXdbK52Li+dSBE9+OxYCe2J10m9cfOMlZG+Jl4DJ1C9WGF9nTiC2OP4KcZ9v9Iva
t/VzWBl/SWMau0sm0d9MVXNVBUkiV17l7MKe654364NSJCS3AJb++7Y5bhMucJTT
tfuenKldoCCnNMrwCrBTCsji1IflrDbPCY+zXTCxNHo+XmTRFSnWVjxnJ8QyAwc/
D6LR5I/PMR9AS7J7aAfF6INeY6qzhM5YEc2YwZSEjoSTwLBGmf9h+xTsVqIavnI0
Ne/bKdvYAq825jPAEV7KrBx3iiRqViRk3ZVIU7GveuzxXFFZRh/3/yj1gKlY3v9A
tihrkeTF7YFZmEOdVsdyQSToU2SvFDc1leumqRiZXuBCpXbePW3kR/VIk5br+2z/
H6py0QG9n13ofX4nw+nP3pgh7XyzL5InpUtu1m2KFy8F7iieZQyWu3EAK0MwZA4O
gz+V7XT/fPQjyP1CkHkrLCUXgUymKziJGyoppJsGMZBbiKL3YN+Jqpvqp8zkx8VD
n8EZNbIksXEuCUikTpipqMf0q9OjFpee0jOvi4JUJLuM+sfmMzh49/WbExFndd4O
cD/qmpMl9FoTuDKhKXOf+oV+qIbzATlq/nMFIPbZxKdcA4kCMI6IZ6CabS75yGez
HZNnncfS9lq9x+OIKipeh7b80PYjuWUBDc2dW607km3b99BapSfb4ntYTcTt5WRe
2KFQ4r2B6URT0gW+cUA7cyruXV54OO5CDUxR9UT59MnZ6UqwV4gbQrboTp9mD86q
w7upbgFs5t66YYWvF4zQGDzXyQy32PYA3wVNGe+ZFF6CbbMgYFuSoynAT8yvvqTY
NIcTymZhXCoPlhSRGNg6RqM5LJNvgx7u4JSS60XdjBEQNEFOpgXn7Q5Ek7JHRo2r
wcjbd5pQu1yb1JRLbVsG9l3MNJ2Tc/Vw5TIRg//9I5HRfe/GVZnNLm1atc6BK2kU
EYJptL9A/timRx4mn1TNAzQbBxBhv0WVW89tTSKdovfb8T7bniPcFOpJT9HAWT2I
AbKAwJlK3XKmKe0eOAdAO4pdZdu83BPZ2bq2a9jfPvMJKhkMwWzH9reG+YzmBKOn
MByMDnFX7UFGJ7ZMCPvahDepzf4g3wM76yZHWbBvRwRUEpsZMIFdAVv4gxf9xwhe
TnR15n8xcLEHPEMVxCjWFj1c82EjSGRI0q0UnHfxv0I+vZqkXhZQHDjdT8TBUBOG
V04B8rxl3JcW/iujMGGHKVIF0ijmL1FB9vp8XWLlVCgJEjXgisZdWeTOWI6AGhhc
cgAiDadqvAC9IfVs1rzD6jcmBhvWD5PaGvMxwaILrHvgFh9HP9z1WXW1MnTCpLaS
cUjRzFu8o+vwSQPtsiJavOAwAi54WvV9dpbQs6HY+OP65kkYyH0G1rb/1MEwW20U
AIWplmAqNfnN+qKFCxdZNYQJH7f+eQ1IJC3TQSATEig/rR9Gms8TgBouiYAeshNt
RwkAkwKk8LWn/J1leghv3Xl3tN7w8WQazKRUgc7PyT30ijcar7b6nga5UMN5zka+
AyGjFN862P0KW6r8VZ3jMd2yqp2scTMu/8smKwwLdq+ncLAstSDrWW5tTmCqr9h9
zS1sBRzlFlRvP+kPpgTITO43Il+fiOLM4JO4TPwvnwz9vgY9F/IhZm9Bx8hduRVg
JmFh5EOKAU2vS5semc5PipukQoiQxjTh8fH+ELDutrZzqF8un4ZVr53r14KSt2oO
g2c3R5JoZl6IZ8yxoH9wRl9m03tgWQofpIuQ5MAExN/LJPovSxgjObB+aNAbLIQ3
WcFgQfBVgXOVUE0AFLM6Npr/34qx8kB5RtoZJC0Snr3slWgwpINB2zRBvEDkiSEL
Q8/IGt1INk9fxHjd8PkSljBOFcAxpDkavJjkKibgSyk8go892/v2pohT6imppE8E
JD2h2To25ciHi4E1wr2Ab2t+V5gFdX2E8rcXAIjNwSTE66qltJ5JS1C9UbEdR6S5
q8FGCFCEn8w6rYtImGT28XUssmmMJiFUy7qiEpsKKSGsqCi0/jw7xhyZPMhO+AOO
lRC9LMNUv5XUZf0MIhxZAfeTmOZS0tTv53pYM+/pMgCHypoFe9KXdRyF/uCu04/b
ho2XxcMpfeGPNGchmxUS2LUaSDDbvnJLnkDqg43xaBhz9K3WKtkHfc4YfAvYh3XF
zZmbtmvUUTjhlmysUepYaKIG9dWS1WJet9tmpVt5Tb/2lSWPUyGdpKUHFeoprBnK
lyzCNXix3as40S/TAibjqth7ckLZBMlIrgamN1pWrbxk2ZZhz0Z2fDS1y+1y2j9P
GfeCkyPsLGzeElqaidAaOBNaDPYtgI7+DVZZXg6ZN3cPZUXQtWD7jymvRo2v5OGn
VHozrNjYIASQEnxO97UKywPZB/Awqv9Dc+jrEzCavHMCR6wqXlR2gOQ5qL3N8tu8
Esk5EdSvYa4oUWkGKTFXdU/MM0tgIeQe0zxpQqOzM0SLL1sPCrh7JPUEyH8BHfK5
y+XJAD68CBnsc/DHXlj85kK52NBPa0D1Wr1NKm3yrwzfMD+sYxA9fEHMrHQXQ/Oj
wUTNa/wBbISbjZfN3l33hCm5bvVVZhANbw8EAWkxrT8GbJ+dXF5xp2NXoOxV7m6E
/uFHNLMb49TEr23igK37gnqzpQKEoW8rpeUgYmDPDi+74naK4DEvumPGg+ppbTgR
fmWeC4a/xmGyYhUCvJDrkn09P9w4jXBBGQ/5JMu7fxypAGSEln6Ntf5fODi0QrRG
1fFHYnn3UGhmPU4ZAs8GKKRSuK/sFYRdwRQxRdjejaYzoORNDtyUJLmN2x7UtM2O
x0S/+li5YTEsZNnnC9FF6rpj8oWmaWM27sVQCj68VxJHev8qYzXKVa2PySp2HsuS
NSLR2jItFXOD459Pjb+tse6/l9vwEo/YbLJc5A1vTbp3JbNvR3et+sVyPfezATJY
0Y9S4QXX3HZem/OoPCgufqkIv3XuMEdxw/jvPo+07yrOim/DNfeCjQxZ23dhK6uT
DR2GmVqJu0L+BuXrYo9YN7DSGyEsyPdX7r+Nx+yhAeZCK/lODKNUYmv+xWkE5wTI
T/lbmtgtu/9iKfFmJYw+Ugd8MIo88ygVKhB8+lQeSMy1nr/v5zRBIKV3vuttywy+
J8gMgl1CORrYI9RGjPjXbdP+7BEgi/2e7MlhJoBN1Ddg1iQRYzuCnhFQlB7pJEVT
7dBpnTleGexbs4zWeg82tm1ZFPe6Fivph0npqB7aNrTnAVjJ5Qk8F3IlnCAQVGlk
7H5osYXzVfbeW+vsDvMUFGXX5KUoVbY8Ot4cS70IhRVLmWK4ZfRshUZNP74NSYkI
NxljGRH+KZ0Y0wCAeuRsVCTzMwmEJUNKOfuzIGvLH/6Uouzw2Oj7lBKGqpD+jaK7
2105wiLc0s+Oha8djSedN5YxvXpKFjr52GwaemS8LewlVO4jmgOc4QZR7oaJYFMm
Yzi0FwHcNmoDIbpSm103Ynws+MGiKmVeH7IFYZgD3hjo0RELzDCL8nfYgHhVofO2
XqnJ5q80CKks2GiHAtA9DHvrNefg9oyR92wQGqGWGxBLF9bWGP5O+SKtePACmjEH
y21vJKxqwGZl+GZsMrxDCRXi/rrjCZSiH0qqykxQiuzAX1eKGf1JqpEM9/asbqtH
S0Jp7free9Gc6U4WLEULXFs8FbCaaaRdh3rj380WnYqwITzjzwMj8ARxB87UPKKO
bsfn30koCD+ok23oy2g7nW995CkUgaISekLJnRiQJuUvLQp2YxG0Xr/1057Yq+gl
OYyBM/jN7p2eVNQB0L/3l8JvAGrtJewNxyES888tgsDMSM6vA3GWZXd4w+VF7PKW
N9OD8Bej5cyRe8CAP+/2UvAiX6rbPT0ENnk0O/GvJ+Sbseqh3x3sm9zQK4qvINzY
V1TIJeIfOanqEASsg0OpZFJaVlhMZ/a91Uc9X9PFhKwjmy6kQT6UZhLLjc9PtWzZ
DhwcRCWSITdy0BymN2hh3PUG4cmPpBeIZbRmqvGdzjZpClhe8FY5tU18tVf0N5VK
SnMptxj/kznywdCW3uCvUrPgI0xBlsfN4rTUhnZ003Pu6qQC/Kn0WRPTWUA3zkN+
mb2G7gZAK+YYoNQTXT/ouX9URvXsPRK7L6dFHAe9SXjynWHhJzdZFYclpYalvW0y
J309jf6GlU61E2wjcq3RjQUykQGThW11PO+OGlpOLhm9hzx9woZb+TPp2Zz+C8gp
CYBy6uYXxLcPLEcuKBKShY8TzFBpS2GECqjoeKUKtU8JDXmkM5z1djrbWeU+wtQV
5/bLFXGm/toIqF4NBQWoMl623ALrnvoDirQ1XO/XKGCf1jP2IdR1pEeldo80f+cM
QS+es30uA5IJmFV3wi4QmB0lna7+mpjtHFRD4pIPQIbosIbw7zSxaO48HvLhz6Ui
Pti0J9EbVIW9HT+rv3BVBCAj9oo64ediLDB3s6jKqARnesE8gQSoB2Gy6tQfzx38
07vQeWFpr8UggmrY72Z6/37ivweJ+xvq4+hs7tU6NNrP5e5cx3Q6M+ZEeatPanwf
ZtECxCgokxukNEvSZUE1v88hHe1KFoYWmz4ODfjAZ1w9YsGMcuRdlVuSdZi3fFIc
3mnYoq8R3Ex14EpvWV5VWxtEcUqDQ1bvxiCoGmHX116lP1ve4u7pBEyK/Jxvywp2
Sv/dgvSOFAJABBcrnZ1vi0HWWoM0YnL47gWeFB7+6rf8SsDIQzDDRgGCb6X6/nrl
PVWyrbutgvlj80rDMMkI+7xqS0hRRftlclBNOfqCF8YrORe5qjMa1Fqy0rNfpK61
ok6kpsB1+uAG1LaPToZ/Q1kOnMJH9Xp0SOGeY7PfH592qChrd9jiUmxpfGUvZmTt
AxeI5WwgTub4GFmU3vEJyJ10wn6YFjca0+kRLi/3yl1ORlAP99wfugEauhRrqagO
UjL2EkOd2c4Y70faJiuhtSaEkPc2HmkTcYjPuM01CBmctUrgHi9Is1jI5fBwHSSL
7BZjiQR9ruc9yZSmNAfRFL/k9XLtZ9U3sZ+kNm7OYIsAB/7ls9dD6tLr0RXab9MN
ceu7w+ci5Zp/8m8ONZco1X7ET1yvUqO+HjPmUtLPM/UI64VPbOoa0KR64So/s5SE
ToKNQjG2n2mSeHZ1VjeMmkN/zdr/5zMvhfndRDjdX/2m8OR7Vue9spSi5A/pRvj4
vpzun7gdK2kg0879zQeCo2sTcjkiVF8y+a7lRn+gcGZDpz0jZ9PgJqPVj6cmM3ZH
D4aycHPUemIRTFRIAgvmoQRWDNpiQrKmP4iehyL5kv3NBohwiqTkd7Dw+j1hGHGn
cEzvsY6XgH/s+uu+G4Em30C0nkFcGGMzq51ehO3S8mPznSZwtwLK+W+I2x9UjI85
RBk5fxN0C7PpYj99BxjRuloSsDdos+kMnhL8t5S8EuMs56/FzPRKIAz/+rqmDQCd
PgLUF6u21W6u1xdDUR9hokyBGclauPjB5FiihQRvhh2VKgbxcpRlE+CDPR8HUPsP
L2+vrPfU2gmWqBreAH5P52FV35SylNL2xSLS31BBW7O+/yu7GiqfIT0BYSHAqJQo
HSEOeRwIOxgReKBXzTMGDXAxojOKOvdwOHdeNfmRLzQaQ5wu3OAOEBgdXjqfogFk
s1FejoXyqtHeKHJEalS3mP8YQCdZWTh1nWNh1g7E7JWBjUpEnEPuk1YhQ0fozkVV
2APhsS9lmdXougIgFn9aqSDMfsQfcYEyzylu/rzVFpUfPiCFK2lFpKFgyyaWu03W
SVsUJvGmiH0e/V713AODYekaKeYXrDjLtjR5nuUb+Ul7FneCzEgAxLQb/wtLyT92
ohbQk5E1KumRocuG31XcVU0UrEj/6ZmCdicW0Yu6WDO8eCq6pYX8EQYszrlyOg/W
CMJ7MnMnGyYWDBFNIyb+ll/lXVs0ogddK98eFmNbIxkdGlvpfn7qsvpzHyBWOvcr
Rj5Q0G8XiQq9PmTYPl/jYLZ2f/RAE2BbZ/7QrVOpaEA59DhfN4g8yiYW5/eUgPNU
SBy8G+YIou3uvRCJMbxQU7d7oQHxyCrnHHbulUaowJ+iPs044qQYoHwxiVlsR97n
Lrw8Z9TQGbJftBrA+04FRsZYaDwSYpBQcEjXFPT45TxMOzlwv/JOVft8fSJbSJ/A
WCtrLagtZELVkjNq3KbniLIwCwJOHcjrdkdul9JgJ+5heqCDGKDXrnM/k2SSjBxJ
GpSciAnHYsbb0828BM4iHR4NFuAZFQS454Rf2gnOYDQ4wxXPOwxT96fHzo062tFU
6eY8Lz8R3UW+g5icMWUzN8IuPQwwAtXxo+2BTkvG20+4PqYCDGOIDGvcWJPlLLOP
efxjNK9QJdbLNLC62pLmAcQoWvWqvKjCcz2Ycy4J4/EPSIJ6Vh8o3JXk+BFtkiJ9
9HNsnEhBaeqphY0ZoEx8VZh0IFYk6aaJ5XrkhyN5BCp0UqR2R2xq4cLxcWM39/9k
k9b3LBGFZFCABN6y7qn6dBtRK0Aad1ddmPG1sl4pQHfLa6rc6KNdZ4Ze1nvZI8O6
folIDW3x6ctfoUB/tvI6VXgFFqMG3B4zY2yN0mMrKB0k7l82v3AhR7nZg0IYOWlt
7IPuK4TddERg0j4rZWJzs6ii3mW2fv62LU0QSPKBoRyAxaVzFzVVsgsVt2HKYlRS
ZWf4SkhMHZyYde3VZrjVcOQ8DLBulAOfV0NsWctd/FGg/MJ/klCNqxSNUGjwxkqN
dUuMmHGC4msCaGrueGVywF0k99OJ06uz51xb47fpwc+wG5OTJJPjLbnVIo2UKXq6
eKjY62QjcKJUtP8KcfnUDajb0A8Vwm9yi8QceVP3Qn05NkR4Cugn/LqcF+pk2wx9
jEM65uTMRM67A+HLaSplY/D+Py6JRXr5FYfPODFkwxQLVWBNi9GQ5lqXl6OjxBQw
t6rwK+hWyyb7pLZcDTJsKD1WIVeroDV9gHPL6Y7Q1fdDXMJfNIHWIid9YiCnZpmT
n+HcquZEjRo/ujK/dhzBJUHZAIeecytYsUlSjIVBcBct5yLk51cRWO/pQx33adD5
2CHfUjj0CVaE4QHVotcmcxzCvemzBtaWLaTtrTOkgWYkdoaSfcT3QVsyNOeDhcnS
pVU+5GuaOVt1QJFAD1Iu5dZepAMij4spAAQIYpWZniBTz8dv7GqtjviIN2PZSOi4
4wN7f8Z1W2tN+UFQovtO2h3iD+KD5zEGmPxCQ7twGuYadAsWiAcu59W2BKLqwjdP
LqA5USu39SxY3DA8blcRX1z+WzM1wQopU+Ye/LzSQalO+tHLtJJ9iHwqVgZs+vVK
5a5yScEPKxzNBaVNEevWjzy0Tb9Qk/aNfHSQKbE4ufrYrc24q4qnPS1YkTBKYpPo
bQqFH0d84YjqaReMEZQSmdW7sm/GOhVVxHnFHyDry4QXSd1dk81oxP4OcSsaA5KC
UvpDcipIyEmP80hi3vy5BoOuZuK3MTljOTyyD9or/wUgtZGYrWlQWgxHy4aKXneP
LrJCHrdW+0WObPV6grLSwte4G5I0BUERNmtCr2O7ra4M/2E8Ayu5rgsBGrJxaJg4
sRISNd9fYdNkpKYN/GBXWZBNLNxwSb5jsaxmsGREuTgwQ5Qc/XN16wY0kO8ouc+k
bDhA9XS5mtY2bpoKVN0vXBrQb7Xkkt3LVifn8/RL/ZMM3myWqZSqUEUCZfSxPcdu
FCSEWuRBdbWYUGXOAx7fK1i0j8NSmtzpqEe+q5BzPL76t/iNaL9TbWGfqGlRioD4
uXWJA4nrzhOnSAEdFW0TeolOk3V9Wo9jNPj/47SguuiQfUKxOxOcaIaZpYpM1mOJ
DQj1br3QHtIug51L0zHcDhGXrdOalaZhZHE+KbMRqtCY8YP0j8RsjlaV0M3Dgldt
WK1rd0GYHxVcLeM6ifdEpApYaNS+TKriav407CBpkyEp9PP7Ujml4KjwUsO9ptkQ
c5hN3PoAewkbrh7o2Piou4kFZ+CQ81OPQebYj5f7e7p5aYRpq9j8Nji7BWLqMUzU
jLHJL79FnGD01mAA5/dPFm7QqyDCUZ5c3uvd42krcP5c/xSFygHLCmyM5RRYdF6H
oR80JozCnljzUtu8FAfj4UXhp4wgBN0fsu3M3Vd6OF1PkNzF8EGr1lHtw12ha+Dd
qu8/9BqmXunj+YG9NkZ907NJ8U8CiFxUeeOj8VHubYb68MaAAhPatEerQYytvuhq
wtWLOqmh5/ZSd2HU/vVKJgNwpxRA4QIKCO5gc3fnOeF86fovTr87El5hinnyqaig
h8a7wIFAMkyuGqiC1CPVX5++NW41lvTV+BgN/QUvWlFxifLicf2FGZ6SCPpC2oyI
jGsFHufqhJmvYuxX+nXnE/Q/5QkCTOHrdBMGxPNWdiKcNBF2Ve/ry+vGiiFVos0p
0U8xw9dKqCeNeZ+0G0D2RDLODDnguHaE2n3CmODkIHyscNJ9yDyU1knQYpt/Tx7Y
jHARh3GvcEnghVnwhM5kklJKYnY/UyxeyvcvddrXULWL8NQokF4fH9d/Ctn9RJDK
LPpmPILWIfO5uFEDg8pLhqCm8hlFTrv6yA/nZCdYsHBTUcTyIsJL8bLl5n76hiKW
1UhnXqHB0Zk3742AdeGqXRPj/a5cokJn/WmMnFByK2Y1lrQjbJweHGcH4XSFTMDu
rZ+OvzLOfrB0MsKDzxGBsWPh1dNLtAAEhlKOdr3/+J4CbPi/VnYich0+RxDq7cHt
0QXzVsf2TT2mm7yZYOcoWz8svyCb9SaL37xp/aRgQ2yRvxljImutuuAxuiCD0A7x
2HYjwvYcZvKZUc6T6/FKa/ZqX00hGXmR6VlEyqIKAT9E4biQJm8/q80IRPoG/kc7
Y06XB3scCDFv2erUVKMtydLRvxeSVTfysFH/01xtfUTdVRaOA3WbZ//spYcWT2CF
iVUwCjUTQRsd7c245SOD9ULxHj3PXxW2/bDx42rA7kTF3ln8y58Y0AfHILn1ykk3
D29ue6sL5C8yCPtoEFBftwGJOBSvDK+EhlbAWxprKZFZlrrJbdVXrnqHyiEpL3qM
RdTOlisTKTaQ8nDIQr0DMnQsG3SWkA7ShUq3QLJOjiVBfvpw9efpQjrY8I1Wc49L
XxBj5XFRrvWIa6Iqc9FmYVuik4coeF4GSLq9nVz1YF2/Qw/gsHsDP7dyB/dT/pRj
6gHvT0IE95JhcrguRcPu1mLHmcEFAlhkXO1jjMn6of6nt0A00ICKgQhCVW5eez4v
3FtkFOso+QyHxGI+vFj81Yb3QzTQNwvG56FlN/AwmvXpJN/AYUGRmnxlZ8TnsppE
VVTRx+1n4JT9n0N7h/C8QVjxNjhpMzMTsxXYIaaeE57FrM3drinYpTvTcrJCuOOu
8rsNLV1x2g2TP7EholhP2pKaK+yByx1MOGP/tbVFv5bCNOPpw3wRPrI7XucIcb72
jvFOpelfu5kImt7garysOP/GpXRs2k1ooDG4Bo0/qnQdUWa5K4PoXft+vRQ92vhU
SyzaR5tPaeeUVd++KjqY2Lr6RbzECVEAMG92Bi1REYxJAUlAb0nmAeIUrps8trsL
Zf+fLpVHdixX0cdVKI+ul4rBMFLuj4u4RCCZk4XQ2q8YPqNBrmbs8MllGWzi7BxF
+8Ea2Bz/sPjuxNUCKqV75c1Ps80yvasrF+35rvbP9ivn2xlXlWNhljtc3TUOajEI
FCVjkZcG0btEhy75k04yFGFWI3ufFmWqSWT1ZhwSzAhUhfkvJf3Mf65hyUpNwIKH
qLRN/LIJjR8gmD+x8zVMQi9FRgoNRM7MDzhccgbkbsH+zIVYtWEFyf8IfFvWRFNz
Job5kFXqY2xGnp7+BqKNiQROwZrUPnmEjXRcv8B/bdDWBBtvsK2StV5LyJeNsmf1
Hw5+VK2q79CCLttaenKkZbDTFN9nDmDLcn2zA/KbcMvQW6wzeluMfFFWNc3Qfdzu
ZlTxh7MyA1gzs/9aLBZWRDI7kpq8YGLydIHRIrBNj76MMBBQH5Wf7MEfADI8icHk
Gju6C4zCh2foaXgjJ0Ws+VsII1VdRZXV9kV9Lt2eDOudfI/CtzabVuPYM+m+bPPD
rG8pkqPeaIFj/v4z00dSZAsbG0iAZ5r1lM9mRZ5Hq8GY/6lDoK4QkGmCkMIJDpnC
eebIr+VJsrhVMvwCBQVAJfNIG1kNB+Yz6AP1bG+F4AzlWo+YDcTNJ/D+Ei6acSRq
tQ5DZ9hzWrl/Xw5VSgqRcURfOskrUR+GI3CvkV0LBK1NFvkNPa9K95Pno2fPu1Cn
kUZwd/lVORNSXZWhDzyhCuFXRSokKol4ELFDB5LcqidXTqdgsOLCiSflqxG1XLQv
1ZzPc2vMmsQze9tpBsEB5ztzvUf93uAiOQP+qjBGlbCmqJs1ls7PWjARDmxYJU61
XeDalmcujhao4Q4VxmCmntONKDZVpy9r2hwPiN0xAtsPY4me++fS2dSGxrlzEzoB
Fa9Ka4IPF3oTkuWTlnI+UetiVgwqDKamNIrA33jByG21c2D8GW/pM1/HrhVUHInz
re7pigxCodbuMcXAX5748Y7Wwm+1rtAV8w7/iFMVfd53JLU6kowdO9KT7MYKEXbA
qYvK2a8Wqc4fFbPIa+6H+WzWznJ2qATWHfYJ6nFeRSTnSIMSi9waiRGUYt1LhAgm
fAkT94D3r/PK+20Wk72Que0bqA+D0ny2JlwwCiGdDKylUbg98tqM8hSQhh4XJpOF
8BCuWwhaUHAv1S/TucYnh7d7OmQ+1omVsPTVP/ftJnVVA0+0lDEug8tx0gXEwpdk
AlazmO4jdXS4BniyPvhRD0z98hBg3KwYmuIvHNfVdrO/9a51jythvO/MrUtDT+77
N1P4PsESc+NVsF8r2IdXienEcSnNXOoh+7CMEJ/LUmRSTKsYigONvYFxF/yfFkRU
LCkJevo5gM/2rGiPNMxiX4xejwthmzikceQnlq8adQCXJMhEB6cM1TVbyquwjU/e
SpiYEBJVI0OxCKax9uXtuzSAh8qDzvsRJn73BjTToKh9yEDKfxZJy1KJWl8O8OO6
K0WuNm8Npeihb4V6sArcYUM3aMe7nsKBH/uncfFjsTTUaBQk8GcViT8giL2R6Moa
DMEnAxwETjCJooZSIAqRIqMLlBEUqTbhk0/qB2YomwnPl0AZEO5+aw4RQUYJlbmy
wfPLh79XzxTyGMFecrQlre54wBvus6enlbFBmny72zJHlw8YEck2rsEtNlujrAph
ZTDZcetz842pRejSvKqfPxPYcE8R1whxwu7NHPKApJNykCV5Kurc/P/A4qu5/1+a
fBYgt9kZinY6xSCtSt/LintEDvCYL4TAXvIUsnsQpBDmLVxk1Pk2bbScboMvHc+W
Kj0gb66hskF7lduhg9hdU2nMGN6kN2wGBFAJ9ntmluX/U1tG6WpDeoLmEnOyBZxx
/DABinsLzvPSwjrjHDJ0ggz7zFXR75/t8vuhx/mRsAGBYqvyBPmTj4dQ8Xz8Fenr
lPMl40HM/X2pVwQI/HFrYc9XmwC0reg8LLbwL59dekUcsr1JOG3HQSXwV6VVmTyN
BfQKbtC6uYPSg0NHkO/ICnHet3wevV4uATBrYwWG3CBTO9eBjSKe9EjrwBvFehmc
GoqfzI6RZmyNzZd18Yv+fnLaiWGNHJZogldKZRIv/RCF2vPJLTtHiLYFNTvlNhbn
8CnIXOH9LGANO0TbOreJD62uNvGBx3MDLvmq+RAlnyjqU6rsIWNakk9PccsusUfy
x0ovda4b96SHut/fjIkJdmL62qYoQR2VP3tZpofxu+cXgO1rx2K2QSg6oboa/CR6
HDvp/e/V9KrYb4n30URSgMrNiOUIcJSGp0rqTzmmrY/bjoBa682Ty2+lQRV+5sI/
kkIVdsT6pWLZCkUEXx3O3Oeeeov623Zp7cl9RDWM5KKW3uV4MwvXiKt04xUsz3XQ
5HqK/a4UzqE8tzdkY6sEoptAMjBgJYsYDHtegcHd8f5x7bT2RxWzWxYLC1qRyaGR
SQnio/LRVotByy2mJjMjdu1FoyLx5zFJsYiC3slNKaizhlWF4vxVby+ZvBNJ82Uv
eq5XD1HjIZcu0dUFrrMKnlMlbYHUjR15pTfyOttXvmeGWnO4ipKbG/Usa6bQnBto
HVrhDa9ClZFqQ0HAdbwdFNQsbB3a10GW+419ZSwRWYDofrmvSifWa7mdIzit6H0z
jrk818jtKgIYr73InrBF8Nov0n2tgmP/NaVjnezUWwOfZJVKTuLOPvjV5qYQ8UcJ
Bxyus0EF5oKNcXiaw4tVtI0NgwFLexiemiQW+LpwSU76exzTlEne9GxJiX1TnIzR
wRXuJK8tri2MeMnWNoPYkEEOWuP1PngZaxXUs9HqcDxXrhWO1/u1PmLJx3jcKH7k
FK6+BecIDe8auS36jWTtUN5uii170QFNAjgNSgF11OIvpRhjfiUvK7H1ktwPrIjf
PBRzAHw+426t+e047gVyhh2RSt4529f1aIfqbJ6XxI0ilpI6JY5PjF2qCpRG3zDs
whI8oJ4cJp20bv/h9LWuHRDzLsCe3GIVopkala5kviPKZwaS4CndHNRYcoa9nmKT
ixNQHyHLXdu9eQHDXZz3tJkmH/p1lS9sTjIMj8VO5G33oNq0VbyMmywrmtfOBTnF
eaKV06RIyi/+t+ZW+e9y+0T8zw2M+SttAF9H9xuc6f0U3GGwv3WXxD1QVu/ZJDbY
KP6PVrhMR7Ht+17WVrpUYbZBfutX1NJxOa+1kBxO+bzGkHZP4/87+V4gFLH/KNyH
LUzl05MqZFLnyA4kfXmPr4dBxvNRQJu1L/pRRYG6Wf2bapoURdv92TxYnLnFr0Xy
HttkTXB39ovnQGv3ERv4SHEPm4110TudvVEqO7XJiqF3BqScbyM4Bo+4YdQsUSxD
+TTRkMyhyMEx3EK3bfMhiOMTLizyMvRYmbdiwipNsPooql1toAXURiZLET+6epPm
fOtfPEKiRnifAPYG7W3GBgqUW3EHNLW/ftLvzs+/LPFP5qea0LF0L9rlDn7A5/9u
E7bHf/VMnb4LsjJFRRjgT2c29UJoKqb6WQoVtW6QyVVQ9usc2Fr1cKG2FZ4qbrTD
NLZ9Bxl3Z0DEhcCGFCAYFS4ODGHtewV7quxiAdiOGn/ecb0dT1ryqHOHQnk7c9dR
EqIFLRuoSaje6hnkb1AyMEC+XpQd7ZDuGYms63G5+Y4L0I10brxaF2ymqlraRL1o
V+AGokVOU+naWldLwgiMVEqcpKU7pV1jFmmked0JXwmHo2ALY/lGrU7LtICfOP20
zSEeXkIesemkgVO11ASi2jqsr0zjfo8Qp2FDRW4Zco4jfTYvtl8IRvmsmcAEYUlR
05pe3X3aC7+Sy4OlNcvetMXw4s0K8KRDm2M2NZ72dStMlEm/Iskrsq0Y3beZ7ZNv
yzfGOvovudxDK0V8/Cw3wVLvmEm/ON/SJhgzVszEv8kKQgJ2+PoJGZCWbA+WBnHz
eGtVbairKmNhuFVPjPAYf5QnzBzlljfwTjmtc38njtP0OYHC7jzGDE23EmFl2JiJ
j29e4E1tVlrjEFCuAIK1Ireb6atxYATD5ShX8purko73bPOl3kGkIH0R34NXS8Mm
WEwLOOVEa8eflEKyjqWIn07bwe33sv7t4RfTNWBNC5Vd0KgIb+4tpuguVtpg0TDJ
zAbhdXYXDyUGpSX9dT5oT8n4zb/rMMtu9TsksMvkjttDlku9ZX4AW16tqA+maQCH
uPZPF93z8zuEKFZy5TjhPZ1l/qiED1eB1QOEPUDzfZ5E/kt99i10H8B8C04xX2MT
3j917QoYjyJTdw/jPAhq8MMxxJAdlb2HqCqlzIizuFf02fooTYh6I024lH5JSiXK
VC9QYl19EimhHJ2xtbIYaqhjofNdjAEMioCQNlzjQFehSx4sv1QD3kpRIedvu1F/
XETWVA5nQk70zhWKspdyIMSj+HXNzSSS0FjCHueeGY2xEuTwo5ORAomwulq/s+Cs
LwdhiUKW8N09bJu62wRMg/58GooM3whf1NR42y3OcDjgN4Scvb++9m57VdVXUxvH
bwPDGM48Cxi406c2wIx2Ca3Kg8xD7lusQv/iHFmyyu589kx6RkiCNlKBpztmHgns
IZRcOsNQpZ6wVpGBq3PxGN7sbwhab0LteNKxMaZq3Z293ETYuNC1j0m4fd2TO2wW
X8jY0fCfg88VH0f2R3rODqlPj/DLOjds51xh5t8JUwh/XIaKKNwh5ENKJRN/b5Vz
HFroccjOpxE6mqvpE4jMxAsRIoeFJ5qNidwyykyLhCkM0INlj+VzrqOAs495M9OH
S/c/pKiEMDgir7FXbORkVTWf3gUDzVCmIqFy8O+paE5FeG7Ck54yAKNtjUb8JqLy
opWcO4XLyU+88/4jRkW93YLQ2HYAqnbcxl0/x2BWYtiScDTmEEvkpOLiVR+W2aRt
/s5pr3Y6M7/+BpE4lJmX9olR0xkPHNKIr75jy42a9SchpE80541OO6AI6e1smLN+
DvTCx1vC7jImrUzXcZ7EEUQT5FZEvztjJ+7QY1EffqA0UFNRYMUUgF+3t6bAreIg
NzEuGkJvYIgqxEtFX+SKls3YuRCHx+/pZizLA/7QpolDV6N8EQXmhA//yNef7f3E
S9sUm9I+rwG6JNc6YkiHAk2D5hRkTSLytMYvZmm3qb09XNGxTxXq6Hu7SNfYsNsz
Yc4TWXDBadnj6m91qX8ORWcNBnxfaw7fP7Lyc5TH7ad+ugqNeJeNLn2tvu8U9UyF
1uWxVEihUXHZbAN3OvRGTr8ipy0Cuh8RZd3VRhBowx5uxTszg1vzFnvLOcbITbqV
cwVwp7c5vZ8Vo0mPXcXu1JYxc9RSL7RRl2HX3rCKa++hK3RNmZTMhrbQXmgm/H40
+tNF0+Ep5jgxtAx3/lbpg1l2f91QpCWYJN3W0lMW5a0qdteGkI/E9NMUW7kjFz2D
Lne3VNdCuqoWWN3bBt8/V/RiqFuvPgMh4sIM+0zXjN44LPQL1grXLrGE5ejsewZC
d4Wdtspr8O/duIFTTWJRLgUeWMt7+lf7QfepVfbwAc9vyAetSCsw4lIM3DEjpYH0
fS0DQ5PWHXVBELcQkxa3YagVCcxjq0fcSIhaMox1/uM7ZhRegNFbKZa40JXl/2AP
roj1NVlsUurldDJkumEGEfR9dddV08ps3UnCYTDPNIvigtO0vnoDtVNsPDnfCZSx
12YLwRjQM2nFV6cMbNkzzJJDloozfuum2heV/h37vImYkvPYQkvq0KX1Z4Eu7qPM
qr4OKTgo2/DHYLfLSo9SzC+a80Y/iSxR7VjtK57wds5zVFEurRAs+cannm/q1I+H
kqR2MLbjNt0ELsM+NvrxJiLqKCrRKEZX4Crr/YccxbJswOortkrvZYTsjRoVzT1z
fLGKw0IOUL/2Y0+mtJjE8W+MdGpWMWJLeGbg+B4MhS3opb8U+ka9LKSrd0bnwUzJ
yKyw7E75Uf6zbnrYTFJtLW1sZBgAUFcPB/f5WdOIoPhw/KOstO2+TkSuYR06Upqo
SVnp/f530QPj4V+q4cfShsUYRU8/UhQbu17ouLzv1VIHZqFfYptZqRc1H2facSGJ
uSUNOPe+CVc0uBaglpwMvhCWGUy1H9dcDeJmVsh9c3P13UwHB/bsmbHouegEtG1o
JMhMxjE/O8JZM8HNBS99uOrEvcVyaayZ61P+nfxHrsNNgvv1uvD7+nGbQ+uzYhzn
fNB3vxGlgpwaC3/W0qkD+bnelAr2+wyE2EP9oaW55GATFwl0GeQWJScE1n2y8FIN
HJIwGkVIkWYkrmE9Zl4OaGuZoPrkUU4oGjwM9E7UTqDxiU36R5hZrbTwcxM/bP4p
sSorqaT5KBitG9G4AfPick/VRdnyFw78UIlNYb2FrrFJ8HCzs8uEgY5iEabqqbvo
N2p48dHG0yodiCQxkX0cll332oGxVOaXKqbobXBrm3ljPeEttV9jwP2hiHiHn059
LCpOZfRaMhU2UbGz78zErjkFP/RNCmtLJaYK8gi3Obc3H4w7iPfikhW5Sy1eo0p5
XYoDpZpyNUQbczQk2ln8783Fei0bsM7AqLH9yfxcJ2RP783GjbriZKmIIFvdGS/M
IZEn28pLovOYn0NBiN2Mu8cGixT6Bi8mrudx0ghoVax3tbFHb88w3lM1nfARsALp
xKj0PTW5WEjo8qGg670NgPbDRkyIFNLcXc+Mi2Y1pW3yeqasGg8DBmq2wxaCb/kD
8YqjFfOytMbFCwO9WJyb1XZq3EgZrVwUGHjn+HPhtVOz8DSqMKfwrfpZhmmav0EA
kHKFNyN3HNxC6KrCGvf1XxoOCkmMaK4rBUlTMNU1962+6ItjrLV5L/fItK1B1zrq
BxN+18uVLWozR7NLN0cTEO0lsrj9DG1HM1YcwBYFMHFq/VvAnDIrNtbjZzhav2a1
zylSZROms9PlQX0hGbloEZis53PTjKkD3iZgCM386PuMuN7/KswrnqxATlRZbQ5Q
8kQ7fnl+3zJmQQN1tTKAvDNl4hVZobtCZL0Yp1E7I+MikBf/jAJy/uDWGUUn6wnA
0EphahrNUduOLQonAIJ8HBDFx0HrXu/DKVy49gw3XZQNQHBIt3bJpFW4Hkam+zU0
nqm3S1aRb47v4eXeghZ4fzYOH8V5O03sOxwB93GUnq9eM1JjIAAe2SD9dhGHf21z
uWG2yr9ClB1XzwJuI2XdvYpQoEJOpdaWeNIzn5i008wIdo/6je1ZhI4OCV4iO6TJ
Yqi5/QVxKhrEfAu0nsPYXYg+xkr/YN16MAw87CNv9OSb2GWBT9gsu5F7nWxYHI/f
5cNBXPMFftRn0/mxjAzQIHz0yh3ThoRcuV/kSRfu7vwFxSireP2Nh7fk6bHT292j
BNhP85cpedfTGL0MSPkB59dqOQ/ksZNAyOwinfniGiArVG7UcjVVqt+K9rEyVBXr
6he5+zZ3O7tfSpmVTSuMZrpk1H3nv6iTOnKymbap+byupFOVdmkzuSYwOIeYx5Ck
cnOsFTCM4bzQA6nzonPirGCxDeRkLf15hVB9usEMsKqV6KFMYEcRJdNXu4VnBsHi
49xTcYBfbdBV8k4u3r/QvZ9mWs2d4rouFIiATodQ+33kyjqxpRBVlO2e7MxjD2WL
MbtCOIhxdatHXXYAAF9Y67puusyG+jF1WYms5rbgEZ70myijC3k52E+qbzGexoIt
PHuMwyhrTnBspkHkZaxqqA6xTpy6UQ74C/A2mWZt0oZ76PwF7QcSIHjFrS3P/w1u
W33a3xWj2kDv89c3VBt+0NOPjR10VFbbF1dWu2rgKRSoMvA5QeVZM9MEAMDJniMi
o+lpNdv+6xDFnauyV1DaxRLSwAXnXQkFoExL00hmPS6PVBktmGWtp+3jdiut4zSb
sGBRMjeyd/lAFNIvUYAgQfEJJBc0ZbvOes4R8ZRds4HdWanqaXJDMkE9q7cdgITh
H2e01eTACa1/2HhiokPXEz2Sinmip5UkdumwakK17hoV/XumXsbZZc7U1Ga9ZOPn
Hp+ZJgp7ckL4UEjj0/DfS6zTlpl/wUZDm8NlEhXKTdYxi3QFudAFfjM/WtBK6aWS
p/QQkZSw1xKAPDyOOY1xqK965WLAVjrXwXawoViqeq2fbPVduxSVLbVkzzUjzezb
T21NdWSeEAyfSlj1AqEy6K21Smj0MIY7HMiYQQZRtfBTXpRAYLtn9e2SyxOY+hgH
MxmOQyU5IAluJ7qYfsBG9yRRg5C0uQsZatjBDqcruuxzwsLLR2B6NGvNU+DlNeLc
C6LQKSYvqQqY4dss8JPS27e1JUOiOLIC6SzCjn8b/tNkhBD1DSwe62LHpjPqwfHy
KuX+Yv48TBDdkfiJ8LLz5D4mhkASSqu7tLSKNxtAh9QdY4VU9IHfaXmR+2x+a7+c
cPMsAZp1K23LMJrjW2f+5TBrMEE0ZalIc61EyFcloGM48Dtz6sruXhRHkwDKZKRN
a+lqCZa+4fMYuaRaI5/LCLJieGoEMs1GrSkKJREi3Z0HSI6QriG8pqy06BCkenI1
lDlOro31vRJhozJiMk303nfKpCpCaClvZDN2rm9dxAOCXp0p0eTm28XHYz3+Kr/S
X+P7qYQDozmRQn+xfWCWH2jntynjm2UM1UMnaLZuZXmUHoa2SYQQjQ435Z1rN+xJ
A8iJFsBfa98wusMxwu3s9ODS/tWhALaZTiDwAVDzDgHkB+qtbQgPPO7AZLiSNklS
xX/pqoH6af7knbylPVGTycNwT70zeLhE46sTu+oZbTyObdG0o2F4AKVg7yfTPz21
rb4UWwwfAKPAiqoEkMKO81angUznilVqS0SgkBIqyLdj/HL/YZ9McdVzrT2DPIjA
3WMYrt9VWsN21/nMBkim/EZCgXqrzIRjo0ipnbRuNy3+cFJHt3GeO0M17MsVl3TV
ywvKO1PrCsmbf2sIR0tsbTCy5eT/xS7+IXK+qlAwL7J6vQDwDGnVEmpG308nsys6
OR4rR1VllosBCbMyZsc2AK1mZYvPk4RPcre0sc7BCRstIMHhHrhjjRGJ1SnwhBiG
mjIwGo9V0zHRFqAYl+OCAd1gRcjo2g/YlqkxPs1Z80JSBPV9AtZioJ1nxrCHt6Gi
FalQBD15cr8ib30dAGC0Tc8y9F58hnGeFH+n1Bo5JJUZuXaqfEFMn3vpbjWSV6vc
mL1bsrTz4Ar7n99P5OjnXzitOnKUdyXIRt8fvLlyt9NJV8+hXM71nuLTUO4jXHg3
oQR+WHZ04iwDc01VO2NjH//iuMctiQWb+6jBl4QxA9ZEGXK4Kt5qmqa3SasAwJFy
ByTJN0QL9cIcTOeowdH2oxkVmaP4BoRjWBZiKPTfMxx5So48GR70raSHdYNB6Sku
ALJ5/kZk2twmQZTMzwxvP79kmR2zLfzyyMCGrhBe0I1eFpzPKkKbz8h9g0I/emFG
B07S3FAUkDF+FTJQuTpV/kKQQrsey2KptnLwAGJMsJad+9MhMa3dU0TIv8PKOO7e
E9foWb0CmKX19G6ntFDYwRYposVxVigsIDUxel6h3bL2dPFriqA6UZBUG8R5TctC
RhuzMr2u9OCqzkwgxx6lR3EimxOhGKzkSTq+GO4yQHFhvdajPO0iYqrdAYE+jhTS
WryJ/vU2WdvPrRGTX5dbA9qM/e1kkJ0E4wbl6OnTO4W/RxfzNkht8cBb8avGgTP1
QTjVmdPJ8qxy7521didnrHYGHjzFDNdWxrQqvx9XmxW1PRCHO4u9b4LKj+4E6NIC
kbIY2B4LgddyC4ME2AbnoXOFZ/yhEkgqq/3gOcLvOQBipYkvFfApttdVWYzj1gHF
fXjnTN4eBdl9qzDn+VAj/pxANjGUWxDA9lzaVuuH+kNMyjHNXTrH1TX2eWFHt/0I
e5yhk8GDr1jkqZty5HvOGx3TkF4IoG8jotqVO0t9MsTtjVtF8DciGH6bsGSjF5Wq
3gK/rOXB3sevz1RA+TQb8Dpfd7HlBOigJDre5zHelz7UX1CU1BNFt/tU8IWu6IyA
g4MSNAzXzAbbGY3tejDzHdnI5HDzPL4cljA1VrtIHBO20HcntZzm+gYFr1YeX983
iuIpjI5RcVc13ZQLXvHmSh3EXQG+W2STJipbuw6zMrvgn/y20vGxf3mMsE+7cmPi
Lw4Yu13H2wB6tZSWtD/Ul4mNQn+/2xpBufIbgPDLM5XLoRfT/qE6xioXrQxxbekl
BmlOyuMUtlOJ15KHX9RvaeuezdlmmfHtngOD0fBvnonAEmi5T7cfLFLOLsJlOhF7
JSHNgAPrhJB3UTyE8OJkAkhf5fhIGhHynzDw6E/TfzqjncV08dRW+3Q6YC/OLJJw
XHgpU9zHmm76ZSsuQV4kPDovL1olCi9w+7hDwm2JvU0TKAjFtI2jx1Bjsh9iY9FA
zHex8yjxuyQkGgNrUHs96IXlPNyEsyslOi+gPf4V7AzHB4ZuDy5WhI/OmU+nd5SF
vcPa6YH9EsFaKZ02SEretMU15h8ztjyZ3meDN999p7BB0Cr7CkmmgRPIIGlmq3Db
6t6fyr7V6eZTym7fh+HhPOjkfbWixOFIxn8Q1SajJIk4IIytoNoycTUXZChZftLL
TuboVrlSVBXon+bYO9eWoxSLjMF6ioYfZaipgpiKQuOiSw+besYqEz0W6YT8t1L6
0+FVyE0bnTMPV8ib38gfcxXoaIBPdVSqokda4QBFOo27O+ZBZ5ZIoxWFWtQZGsRj
OtFdOMc0jnOLbbEtil2V3/1KYmOUcvHqh1OZeMdH7PphKcTzSfDHCiu/cwJ105YP
DyhpWh+ZXlrASvTqxoMzLD/bfAaj0BMbVgYRBo/tChpFYZaVFG712+SMh0Yi5TZi
SBomCo+e4fnMPrebV7xtdmkjK7xu79VKF75/j8ELrhCxRPQGEIdbqVnNBL4oyPkX
6AuwYuRGYCTZy5biurvUYlTCAtg7ijQ4MTUNTXouQZSBAQuU2htUIcDbuB//U4Cs
lae8uDQbeJuITrop6AEphq8QLfm99i+1/89lYcONliQdU/IevwewVkTys85xCWr5
PyinJVZSRH92gcBzQMm79uMWVLCHPuR+xijITij7fuZI7DKWqiBsuGipM9BmpENn
9rnPHnjQJPimqlsPXldxYh6QpnNARb2cvtIw6VtBhikqN98Si77gT6s/6wPqH/kL
pny7OKKH1DYwgUmAnkYne/y9UU/4LyzrfoRbsReqyeXKAdXhdg89buAN+Fki6St8
Ebp68yNGDJhW8s8ud0HqtJbIA9mK5W9qfg9BFBs8GXW5Pnjv5Z6kKXM6CBsaK4YF
YMpqHlrQGVe/i+oF5HPlkOkWWHyGCJ6DtuBjWTBDWkP4ntIpbWSf52ZehA+EiPpS
mzIkoDa9PnIZ2aw767m6gDSC09Po9YW5FFF6yijyfUit6sP71zI1LYnd4yDmgwih
Yq40HO81YiS37+dtqyxpJ4LscnKi3NPVNMaFVjoC4vqDiYO6oMpF3+KKhhHJk/Rg
FM816kZTpmaEaE9V1PcUWId6S2vGqPlzp72XTureMmF588uDaBh6WFgEFDFaHJzg
xniAfk5y5xwuqeVr7TUcT5uRV0eA8FYPTXixnltsR7jmn/qXdkHG/iq9VnWNVRbf
xbJAwFeYkIMFL2x+bZ2na0Lf+2dRycZyQjSBTqdIlgLqNJ/bYwVi//X5L1X+TTzf
e5AYFynXIL3Ry2+xkf6asNIJK2DYzzMdAvEF+aAsn8ph4sXuENs0ZUUNWTJmtM/k
NZAF/pC77WikSWFWI/8M3pCmfnHTO+TFV7CuxXvmBVZQAm/aCw9Ydx5m4eSNT3zQ
0/HMgn3Dc2BS8kqhZ1WgD666zf42KEgbx3AkB8Fo1X+ENz+Tt+0t9iKb3HEZG7cM
Jinq4m13FbbbaQrvMnIU32ePYhh6btKy6Wa1GafSprm8sLFpeiu9eIn6kUc0lhmZ
wNGYvMiHBmc7boe5BDKIUbxezL92JdQAvOHtQQEax6yvmTzSZsA17wzu4zO11Vo6
pazawJRobV58fgysdIfVTPcHgRAgXoYRtJikjtv5qQyU/yYBkGIC+cqZF25R/oKN
DpZr4b8WPOrec9dg1+GbMh+NXg7KjUaxC6zIHpNq4ixechgk3G4WlHnSLJLg87G/
DzaqkmZQ/oxL+Q1ZbZ5Gfsxe5Ekud6U695Uq5KL4aF8ZpJvg/b8hMYlotoQHtCSC
8rlY9j1/E71hYr2H0JcKEV65aAtViaFlkagVGt0A1nHqfclx9EwL24XGNWL3YKlU
N03Hd1xdnjXd/OMlbNfEaf2/EdXQzohIE6HUl7eHKHyDtjia4hGNWvaesyetWkAA
CdZSjg6RRwsXaVMXB5aL1LDbDw7JVX5ov9gIxAol6aHZiVIiLIDGabXr3ZsDgNq0
rHSYzXguRslnQ8iYLy2ESLdM0XnNFz5OL+u4GB2jJrtjFHr2qCT1/QNyCefoe+fo
DMMXIf2j0GnfcQSlJ8JoZdiykRKPqqeT65jA1XixBXO/x0eGrCbNTlfuSg1EDu+Z
aEJvesAh0mtmtkpC4vzOb1vYyo7q0ntxp0C3GHGquBuMeY9HqLYxnrtpf0OP1Fff
wlJcf9vA7Y3VMFTkwIKm/5nTZQUCKwqtpJeHdHKym678s1kZUY9cAvNKOxSS3p6Y
jdlQHFcs+hmLSeOSqXhhTEFzkzy39FrJ7Wi1PrRWa1IfNjjsyXhd30A4+gTo5Glc
ltEGJ0OfgugeOWc8EeIFiEjc9Jco7rREfw078dnsp5IPQc0rsitZ+hCfUOUf2EUd
WlKq5FOa6A9iX4UXGPbTsb5mOkYM8gFqMSMI/jOBIg17kPlFo0h03mOVer/hWax3
fZvZHeBUY9hfV0q4g/lXlMj4F3gzzqDjZdyL8AZfDoucbrcFXKxBGcg57sXeGnrK
J/+Ht8GBa5TEwYomCZLPQZKZ+4bzMa36qreEllPotw8MhDXTtRh90j00OVEqQZwL
1vl1kg59v9XdEO/S9k0Va9SN6c0SnU4xyHXZMVOZULP5UUm1yDmnmHejE/ILcYes
gy81dZ/KNxq73tjzk02ynxoUGl5p6Dlr1bj83lMRZcxW7LofQ9OZI9nTfVoG3IIv
gEG+PwPSQjbtEvHzqYqtLw3zyctpQa+4odyB2bdgngwpQG79x2D0Cj6b0rPeiZgM
6gnr3BvTPgpQBSujIJ3XN+QVlv7ZdOnXYBht2YIgJ5CWBumJsnYS7SSL34KlR8M1
o9d4zUoDu11X0ZtxIIJ4PhoaTmA2rFLsPon9am+gdULlpVs0Zet5oVhX1PhXMkRU
uZwZQ0ryOXCOiICTJ3jakW1z2g0e1zCcgS6c8WoJAmD4SBtBRMEdF3r5LfPUtZ8u
4N+cwbuikfXj3VG2UWgBAOdMWdfHVgyJD4HD5ShEtgsjIi0hnR1xDXD9hkPbznAn
QWblq5srMvFwxFcdKmeOADbPbrXsJ7HGRW99Oxq8HMBVQTuJ39j7N3LbRS7v5Ovi
0dz7/mOJZJb0aGciiIfIaBivlOdEcD5d+IhYIPR5K64/r0sNr5mRtC923udEpbt2
JcLvdBtV3nfyvIsiSg8sNT7QLBNYBTzrA2j51kscJrt0Nra2DMIcuPwUjfK4Kghe
A7qce5jrL2rIVWRPxHbZZ/ZlBuqz6NVjV05kyNV4vY5X7VJ/CFpb4fQC9ypjUQWB
jOHQ8zQzn/QkcRmRUpvjFEstFsU+h1sCfw5/JS3kh1xAoCSWOePr1q4sBh4RnJip
f6HVo0U9inFusJer3xqiKdzkqaiXhDvyz8mnU7nxs0ydhCbXK1qIb7anOskLVJkR
IrdYdMnNTKhEcUH+dff61rD7pb86fHLIzxhDIN1FlfNeoNIkkVrge9Wj1x9R4rk6
zcDe3EsV97gIYX8hWueuXeWSDUjRgKo11U0ehHOd+mxYQpwlk51QjKb5Kubrmyk0
1hXRu6QcCNAEM+DxQOeVJBf3sDr8F/XB9Lw4omaltNbfMReW98kW+wyuDMhelVXF
zA66D0SWoYFYkR8Tbl2OIrlYf7Qt1l0l3Pp26S+HRwt2gUI9kbC5NIjbI3XtSdCg
D6f9NKC81Iui9m1XLDAmC22qUKM0K3OYev/32o2T97jQBJfnvaA4SViIsFphIL7w
WwDDdBchOC4+n/VCPLmP/XEWFFaYoXwm8p0bZt8BD68qSy66Hlfd8zrGdcL53uCd
SuqCp9O4/K3azUKDKe2QmdfWMdRPwytTA3ks0jasrPFg/AMKRFD2yCvPqPX8lAik
ceH+lVyJFneewfpy0uCnmkfSvLM5yEXbZo3pTLlukWr1gm11mdMyr4jYkMIEtfFy
2TtylZiCySi+QopJi9EcDxak5DFVP9RcGwW1we5WGVsyzJjw3Uh6RQB3fGsIr4Ke
8yDpBlIB9YvIldSgzuJI9AEoZHFWeb2qArfQs4jLOjRiWkD0+8ktcuaTr/z+J+Rh
fjrLXIc3YtPNKQ1Q6GRzJ9HCsWnOaBMI3VzzR2640QahKbMgcnYqCpTZvkG7W9dc
c0VyqCwz4uwjYeQtcNHaoYktTJeWNooC1wDoewNGZ+ZTXF94w4JKeKIcDKrWN8qC
plZ5Q0bW7Ry6M+AfHmQpJ5XVToKcECvNgAhBacmh025CZZVyk5HauB7NBr7JlCTS
FydhSqRb5OZzBNt2buFrlPw/ZZVYV8tWbHcR21Xg+7ieNs4//s48jRYPV+nbWxxT
EN/jU4PlDNKEVPsvreLVDIbLpdGxeBuez/DoPQXhFZY0GQ7EdGrUQSIm4bjpwkWB
QdSCBZIdHT5MZSTvWRrJ1RxXkbLyosrv4oGEzg/wzC5ys4LPUN/TC+PRXqZNTs0b
Myu/awDUSHw2k69YPLiMue+TSbse+L2sOxLT+hv4ZeU6IHgKa5c7OVJvqxI9KgFW
I+haOTPbjl+ExHSc1k5nmD9iU8YbLHelhN/heh3VMNBAftO+375el4jduQbUHvCI
mjZMOkhF/v6X5jnK5rfearqubpZuqtSsu0SDPnCXOfgvhaNDBGOaN+baRNzY6BdZ
6J6DJ8x+93fuGiVrLQiPvtaDnlO6TB1F2IwOJl00K3SErfSYYZ3uXc6YM1Vv34V9
v85VeaoCisray3p3TlcvotazWyZ6gpdRgAJSpurE+kC9nP2YtxqZ+Jg1IY/0Yadk
5yDSdLUcHVq3lsZOcJIYtNA8ABi0m8RpSKROFnI31rTO1kjgz6QSwES7XlAxma5W
2osA12Eg8HacDAHQlrrT7IMYwmzadFKRKCNCyYlTiwt9cy/VLpcwk3VnDPMaDXp4
Uxc627SgKuuLdsSTO4WuI0ek2vK5bkcDvqG2aapPoofySEmmTARX0NtqhfbpnYaK
8ZjhlttG5n4mhs40AcGBIo37P8nJUTAq83Uv6mLX8zWCf1AXWuvwfDVjz0ixfmY5
sSvSh+OQYsCFdffvp+cditWuG3A8QoemYfD+5bn25qgQDBTibCbk8J4wsIk8Bhtx
C4iivy8v2OTUnT9eaMsZxkWxoaZLGQZp5cLlnQOjRWwepTsesQIvV/hHKut7PYXH
9+Wl0lX5jotFKcgI+ZNZMNBQOwXg+SZ6+A/d/I31G2w0fG3wCa0TVbOrRV0EF95/
vL/HDR0QAg9tLdDTb/i5Y4M7K6Fl7U/MQU59lykf1//6MIB+mfxW5jY3j/+lza3A
NYO9nsKIljtoHyO8ijBO7pCxpMcN8uGEcQm/f5BXnzmwz2NFWERtKMeTNWbRx24N
AXzwMirjyuOLkbHfdIVL1PZ5BUXh73Kb5lsPyVZ4cE/vD2Ks0JkyN+NQlQEHtQD4
jwP5W+aj2JXxyWp6kpCxHtB9AyPtamZeojsLXgb3mH8kDNL4i9z4WcCBtSb/EvGC
GnWCn8mVmNElna1mmrVQ/TudTSu3LwGczp3dTJVZLxLYSL8S0sccVmv82nOI7ahM
a4uSoaY36B9SOPuVv7u2sg==
`pragma protect end_protected

